// Library - io, Cell - PDUW08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 17:52:32 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module PDUW08DGZ ( C, PAD, I, OEN, REN );
output  C;

inout  PAD;

input  I, OEN, REN;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_core_sa_comp_top, View - schematic
// LAST TIME SAVED: Jan 21 17:21:37 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa_comp_top ( sa_out, in_div, in_ref, saen_25 );
output  sa_out;

input  in_div, in_ref, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I85 ( .IN(saen_25), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(sa_out_b_25), .OUT(net051), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net038), .OUT(sa_out), .P(vdd_), .Pb(vdd_), .G(gnd_),
     .Gb(gnd_));
nand2_25 I80 ( .G(gnd_), .Pb(vdd_), .A(net051), .Y(net038), .P(vdd_),
     .B(saen_25), .Gb(gnd_));
nand2_25 I96 ( .G(gnd_), .Pb(vddp_), .A(out_div2), .Y(sa_out_b_25),
     .P(vddp_), .B(saen_25), .Gb(gnd_));
ml_core_sa_comp Icore_sa_comp0 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp Icore_sa_comp1 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref2), .in_div(in_div2),
     .out_ref(net73), .out_div(out_div2));
nch_25  M0 ( .D(net039), .B(gnd_), .G(saen_25), .S(gnd_));
pch_25  M43 ( .D(sa_bias), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M4_4_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_3_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_2_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_1_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
rppolywo_m  R0 ( .MINUS(net039), .PLUS(net45), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net45), .PLUS(sa_bias), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa, View - schematic
// LAST TIME SAVED: Sep 12 16:00:47 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa ( nv_dataout, blsa, vpxa, dec_ok_25, dec_trim,
     fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, tm_testdec_wr );
output  nv_dataout;

inout  blsa, vpxa;

input  dec_ok_25, fsm_rst_b, fsm_sample, fsm_tm_testdec, saen_25,
     saen_b_vpxa, testdec_en_b_25, tm_testdec_wr;

input [4:1]  sa_pgate_vpxa;
input [4:1]  sa_ngate_25;
input [7:5]  dec_trim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_core_sa_resbot_m2 res_bot_ref_m2 ( .div_2r(dec_ref_2r),
     .div_3r(net0155), .bl_out(net0181), .nwell(nwell),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .bl_in(blsa_ref));
nch  M1 ( .D(net0173), .B(GND_), .G(testdec_b), .S(net0269));
nch  M27 ( .D(net0103), .B(GND_), .G(vdd_tieh), .S(blsa_ref));
vdd_tielow I204 ( .gnd_tiel(gnnd_tlow));
inv_25 I38 ( .IN(testdec_en_b_25), .OUT(dec_gate_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I222 ( .IN(dec_ok_25), .OUT(net0114), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I224 ( .IN(net0114), .OUT(net098), .P(vdd_), .Pb(vdd_),
     .G(gnd_), .Gb(gnd_));
nor2_hvt I214 ( .B(high_res_b), .Y(net0132), .A(testdec));
mux2_hvt I206 ( .in1(blsa), .in0(dec_in_3r), .out(in_div),
     .sel(testdec_b));
mux2_hvt I207 ( .in1(dec_ref_2r), .in0(dec_ref_2r), .out(in_ref),
     .sel(testdec_b));
mux2_hvt I219 ( .in1(net098), .in0(sa_out), .out(net0191),
     .sel(tm_testdec_wr));
rppolywo_m  R3 ( .MINUS(net0115), .PLUS(net0112), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net0169), .PLUS(net0115), .BULK(gnd_));
ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 ( .gwl_b_gnden_25(vdd_tieh),
     .gwl_b_sup_25(vpxa), .gwl_b_25(saen_b_vpxa),
     .gwl_gnd_25(gwl_gnd_25_ref));
inv_hvt I208 ( .A(fsm_tm_testdec), .Y(testdec_b));
inv_hvt I220 ( .A(testdec_b), .Y(testdec));
inv_hvt I213 ( .A(net0132), .Y(net0120));
inv_hvt I215 ( .A(fsm_rst_b), .Y(net131));
inv_hvt I136 ( .A(rd_out_b), .Y(nv_dataout));
nor3_hvt I102 ( .B(dec_trim[6]), .Y(high_res_b), .A(dec_trim[5]),
     .C(dec_trim[7]));
vddp_tiehigh I169 ( .vddp_tieh(vddp_tieh));
vdd_tiehigh I117_2_ ( .vdd_tieh(nwell));
vdd_tiehigh I117_1_ ( .vdd_tieh(nwell));
vdd_tiehigh I117_0_ ( .vdd_tieh(nwell));
vdd_tiehigh I168 ( .vdd_tieh(vdd_tieh));
ml_core_sa_refres Irefres ( .nwell(wp_ref),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .wp_ref(wp_ref), .bot(net0173));
ml_core_sa_resbot res_bot_sen ( .div_2r(net0228), .div_3r(dec_in_3r),
     .bl_out(net0112), .nwell(nwell),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .bl_in(blsa));
ml_rock_lwldrv_wp Irock_lwldrv_wp ( .gwl_gnd_25(gwl_gnd_25_ref),
     .s_b_hv(vddp_tieh), .gwp_hv(vddp_tieh), .gwl_b_25(gnnd_tlow),
     .ngate_25(vpxa), .s_b_25(vpxa), .wp(wp_ref));
sbtlibn65lp_ml_dff_schematic I132 ( .R(net131), .D(net0191),
     .CLK(fsm_sample), .QN(rd_out_b), .Q(net135));
ml_core_sa_comp_top Icore_sa_comp_top ( .saen_25(saen_25),
     .in_ref(in_ref), .in_div(in_div), .sa_out(sa_out));
nch_hvt  M48 ( .D(net0169), .B(GND_), .G(vdd_tieh), .S(gnd_));
nch_hvt  M46 ( .D(net0112), .B(GND_), .G(net0120), .S(gnd_));
nch_hvt  M45 ( .D(net0181), .B(GND_), .G(vdd_tieh), .S(gnd_));
nch_hvt  M47 ( .D(net0115), .B(GND_), .G(dec_trim[5]), .S(gnd_));
nch_hvt  M14 ( .D(net184), .B(GND_), .G(vdd_tieh), .S(net0103));
nch_hvt  M16 ( .D(net208), .B(GND_), .G(vdd_tieh), .S(net184));
nch_25  M21 ( .D(blsa_ref), .B(GND_), .G(saen_b_vpxa), .S(gnd_));
nch_25  M23 ( .D(vdd_), .B(gnd_), .G(dec_gate_25), .S(net0269));
nch_25  M25 ( .D(net0269), .B(GND_), .G(vddp_tieh), .S(net208));

endmodule
// Library - NVCM, Cell - ml_core_sa_top, View - schematic
// LAST TIME SAVED: Apr 18 11:05:06 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa_top ( nv_dataout, bl_out, bl_pgm_glb, vpxa,
     dec_ok_25, dec_trim, fsm_rst_b, fsm_sample, fsm_tm_testdec,
     sa_bl_to_blsa, sa_bl_to_pgm_glb, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, tm_dma, tm_testdec_wr );
output  nv_dataout;

inout  bl_out, bl_pgm_glb, vpxa;

input  dec_ok_25, fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, saen_25, saen_b_vpxa, testdec_en_b_25, tm_dma,
     tm_testdec_wr;

input [7:5]  dec_trim;
input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M27 ( .D(bl_out), .B(GND_), .G(net81), .S(net71));
inv_hvt I108 ( .A(net063), .Y(net061));
inv_hvt I131 ( .A(tm_dma), .Y(net063));
inv_hvt I101 ( .A(net69), .Y(net77));
inv_hvt I102 ( .A(sa_bl_to_pgm_glb), .Y(net69));
inv_hvt I167 ( .A(sa_bl_to_blsa), .Y(net73));
inv_hvt I96 ( .A(net73), .Y(net81));
pch_hvt  M1 ( .D(bl_pgm_glb), .B(VDD_), .G(net69), .S(bl_out));
pch_hvt  M11 ( .D(VDD_), .B(VDD_), .G(net73), .S(VDD_));
nch_hvt  M2 ( .D(bl_out), .B(GND_), .G(net77), .S(bl_pgm_glb));
nch_hvt  M4 ( .D(net71), .B(GND_), .G(net061), .S(gnd_));
ml_core_sa Iml_core_sa ( .tm_testdec_wr(tm_testdec_wr),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_tm_testdec(fsm_tm_testdec), .dec_ok_25(dec_ok_25),
     .saen_b_vpxa(saen_b_vpxa), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .dec_trim(dec_trim[7:5]),
     .nv_dataout(nv_dataout), .vpxa(vpxa), .blsa(net71));

endmodule
// Library - NVCM, Cell - ml_s_b_hv_sw, View - schematic
// LAST TIME SAVED: May 16 11:29:12 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_s_b_hv_sw ( sbout_hv, ssup_hv, sbout_gnd_25, sbout_high_25,
     vddp_tieh );
inout  sbout_hv, ssup_hv;

input  sbout_gnd_25, sbout_high_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I114 ( .IN(sbout_high_25), .OUT(net62), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nch_25  M23 ( .D(sbout_hv), .B(GND_), .G(vddp_tieh), .S(net34));
nch_25  M7 ( .D(net34), .B(GND_), .G(sbout_gnd_25), .S(gnd_));
pch_25  M5 ( .D(net46), .B(ssup_hv), .G(sbout_hv_b), .S(ssup_hv));
pch_25  M14 ( .D(sbout_hv), .B(net46), .G(sbout_gnd_25), .S(net46));
ml_hv_ls_inv Iml_hv_ls_inv_vppt ( .vddp_tieh(vddp_tieh),
     .sel_b_25(net62), .sel_25(sbout_high_25), .out_b_hv(sbout_hv_b),
     .in_hv(ssup_hv));

endmodule
// Library - NVCM, Cell - ml_wp_ctrl, View - schematic
// LAST TIME SAVED: Mar  9 16:06:25 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_wp_ctrl ( s_b_25, s_b_hv, sb25sup_25, sbhvsup_hv,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25 );
inout  sb25sup_25, sbhvsup_hv;


inout [3:0]  s_b_25;
inout [3:0]  s_b_hv;

input [3:0]  sbhv_high_25;
input [3:0]  sb25_gnd_25;
input [3:0]  sbhv_gnd_25;
input [3:0]  sb25_high_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I21_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_0_ ( .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_25_sw_3_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[3]),
     .sbout_hv(s_b_25[3]), .sbout_high_25(sb25_high_25[3]));
ml_s_b_hv_sw Iml_s_b_25_sw_2_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[2]),
     .sbout_hv(s_b_25[2]), .sbout_high_25(sb25_high_25[2]));
ml_s_b_hv_sw Iml_s_b_25_sw_1_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[1]),
     .sbout_hv(s_b_25[1]), .sbout_high_25(sb25_high_25[1]));
ml_s_b_hv_sw Iml_s_b_25_sw_0_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[0]),
     .sbout_hv(s_b_25[0]), .sbout_high_25(sb25_high_25[0]));
ml_s_b_hv_sw Iml_s_b_hv_sw_3_ ( .sbout_high_25(sbhv_high_25[3]),
     .sbout_hv(s_b_hv[3]), .sbout_gnd_25(sbhv_gnd_25[3]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_2_ ( .sbout_high_25(sbhv_high_25[2]),
     .sbout_hv(s_b_hv[2]), .sbout_gnd_25(sbhv_gnd_25[2]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_1_ ( .sbout_high_25(sbhv_high_25[1]),
     .sbout_hv(s_b_hv[1]), .sbout_gnd_25(sbhv_gnd_25[1]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_0_ ( .sbout_high_25(sbhv_high_25[0]),
     .sbout_hv(s_b_hv[0]), .sbout_gnd_25(sbhv_gnd_25[0]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_sup_25, View - schematic
// LAST TIME SAVED: Dec 18 17:40:05 2007
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module oai21x2_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
nch_25  M6 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
nch_25  M7 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));
pch_25  M4 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
pch_25  M0 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));
pch_25  M5 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yptest, View - schematic
// LAST TIME SAVED: Feb 26 14:41:48 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yptest ( yp_test_25, yp_test_b_25, yp_test,
     yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25, ysup_25 );
output  yp_test_25, yp_test_b_25;

input  yp_test, yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25,
     ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



oai21x2_sup_25 I180 ( .A1(yp_test_b_low_ysup_25), .Y(yp_test_b_25),
     .A0(net37), .B0(yp_test_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(yp_test), .sup(ysup_25),
     .out_vddio_b(net028), .out_vddio(net37), .in_b(net40));
inv_hvt I181 ( .A(yp_test), .Y(net40));
inv_25 I182 ( .IN(net028), .OUT(yp_test_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yp3, View - schematic
// LAST TIME SAVED: Feb 26 14:41:31 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp3 ( yp3_25, yp3_b_25, yp3_b_high_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, ysup_25 );
output  yp3_25, yp3_b_25;

input  yp3_b_high_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I201 ( .A(yp3_sel), .Y(net075));
inv_hvt I101 ( .A(net075), .Y(net070));
oai21x2_sup_25 I202 ( .A1(yp3_b_low_ysup_25), .Y(yp3_b_25),
     .A0(net069), .B0(yp3_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(net070), .sup(ysup_25),
     .out_vddio_b(yp3_25_b), .out_vddio(net069), .in_b(net075));
inv_25 I204 ( .IN(yp3_25_b), .OUT(yp3_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yp21, View - schematic
// LAST TIME SAVED: Feb 26 14:41:20 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp21 ( yp21, yp21_b_25, yp21_b_low_b, yp21_sel,
     ysup_25 );
output  yp21, yp21_b_25;

input  yp21_b_low_b, yp21_sel, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I206 ( .A(yp21_sel_b), .Y(net50), .B(yp21_b_low_b));
inv_hvt I207 ( .A(net50), .Y(net68));
inv_hvt I208 ( .A(yp21_sel), .Y(yp21_sel_b));
inv_hvt I209 ( .A(yp21_sel_b), .Y(yp21));
ml_ls_vdd25_nor2 I194 ( .in(net68), .sup(ysup_25),
     .out_vddio_b(yp21_b_25_b), .out_vddio(net72), .in_b(net50));
inv_25 I213 ( .IN(yp21_b_25_b), .OUT(yp21_b_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl, View - schematic
// LAST TIME SAVED: May  4 14:26:38 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_ctrl ( yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25,
     yp_test_25, yp_test_b_25, vblinhi_pgm_25, en_blinhi_pgm_b,
     en_blinhi_pgm_b_ysup_25, yp1_b_low_b, yp1_sel, yp2_b_low_b,
     yp2_sel, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, yp_test, yp_test_b_high_b,
     yp_test_b_low_b, ysup_25 );

inout  vblinhi_pgm_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b,
     yp2_b_low_b, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp_test_b_high_b, yp_test_b_low_b, ysup_25;

output [1:0]  yp_test_b_25;
output [5:0]  yp1;
output [5:0]  yp1_b_25;
output [7:0]  yp3_b_25;
output [7:0]  yp2_b_25;
output [7:0]  yp2;
output [7:0]  yp3_25;
output [1:0]  yp_test_25;

input [5:0]  yp1_sel;
input [7:0]  yp2_sel;
input [1:0]  yp_test;
input [7:0]  yp3_sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_1_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1]), .yp_test(yp_test[1]),
     .yp_test_25(yp_test_25[1]));
ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_0_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[0]), .yp_test(yp_test[0]),
     .yp_test_25(yp_test_25[0]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_7_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[7]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[7]), .yp3_25(yp3_25[7]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_6_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[6]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[6]), .yp3_25(yp3_25[6]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_5_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[5]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[5]), .yp3_25(yp3_25[5]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_4_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[4]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[4]), .yp3_25(yp3_25[4]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_3_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[3]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[3]), .yp3_25(yp3_25[3]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_2_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[2]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[2]), .yp3_25(yp3_25[2]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_1_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[1]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[1]), .yp3_25(yp3_25[1]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_0_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[0]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[0]), .yp3_25(yp3_25[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_7_ ( .yp21_sel(yp2_sel[7]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[7]), .yp21(yp2[7]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_6_ ( .yp21_sel(yp2_sel[6]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[6]), .yp21(yp2[6]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_5_ ( .yp21_sel(yp2_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[5]), .yp21(yp2[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_4_ ( .yp21_sel(yp2_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[4]), .yp21(yp2[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_3_ ( .yp21_sel(yp2_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[3]), .yp21(yp2[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_2_ ( .yp21_sel(yp2_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[2]), .yp21(yp2[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_1_ ( .yp21_sel(yp2_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[1]), .yp21(yp2[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_0_ ( .yp21_sel(yp2_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[0]), .yp21(yp2[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_5_ ( .yp21_sel(yp1_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[5]), .yp21(yp1[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_4_ ( .yp21_sel(yp1_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[4]), .yp21(yp1[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_3_ ( .yp21_sel(yp1_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[3]), .yp21(yp1[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_2_ ( .yp21_sel(yp1_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[2]), .yp21(yp1[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_1_ ( .yp21_sel(yp1_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[1]), .yp21(yp1[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_0_ ( .yp21_sel(yp1_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[0]), .yp21(yp1[0]));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - io, Cell - rgtbank_1k_july16, View - schematic
// LAST TIME SAVED: Jul 21 09:26:20 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module rgtbank_1k_july16 ( Tdo, in, tck_int, tdi_int, tms_int,
     trstb_int, pad, TRSTb, Tck, Tdi, Tms, oen, out, ren, tdo_en,
     tdo_int );
output  Tdo, tck_int, tdi_int, tms_int, trstb_int;


input  TRSTb, Tck, Tdi, Tms, tdo_en, tdo_int;

output [20:0]  in;

inout [20:0]  pad;

input [20:0]  out;
input [20:0]  ren;
input [20:0]  oen;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



PDUW08DGZ I63_7_ ( .PAD(pad[7]), .C(in[7]), .OEN(oen[7]), .I(out[7]),
     .REN(ren[7]));
PDUW08DGZ I63_6_ ( .PAD(pad[6]), .C(in[6]), .OEN(oen[6]), .I(out[6]),
     .REN(ren[6]));
PDUW08DGZ I61_3_ ( .PAD(pad[3]), .C(in[3]), .OEN(oen[3]), .I(out[3]),
     .REN(ren[3]));
PDUW08DGZ I61_2_ ( .PAD(pad[2]), .C(in[2]), .OEN(oen[2]), .I(out[2]),
     .REN(ren[2]));
PDUW08DGZ I61_1_ ( .PAD(pad[1]), .C(in[1]), .OEN(oen[1]), .I(out[1]),
     .REN(ren[1]));
PDUW08DGZ I61_0_ ( .PAD(pad[0]), .C(in[0]), .OEN(oen[0]), .I(out[0]),
     .REN(ren[0]));
PDUW08DGZ I94_5_ ( .PAD(pad[5]), .C(in[5]), .OEN(oen[5]), .I(out[5]),
     .REN(ren[5]));
PDUW08DGZ I94_4_ ( .PAD(pad[4]), .C(in[4]), .OEN(oen[4]), .I(out[4]),
     .REN(ren[4]));
PDUW08DGZ I86_20_ ( .PAD(pad[20]), .C(in[20]), .OEN(oen[20]),
     .I(out[20]), .REN(ren[20]));
PDUW08DGZ I86_19_ ( .PAD(pad[19]), .C(in[19]), .OEN(oen[19]),
     .I(out[19]), .REN(ren[19]));
PDUW08DGZ I86_18_ ( .PAD(pad[18]), .C(in[18]), .OEN(oen[18]),
     .I(out[18]), .REN(ren[18]));
PDUW08DGZ I86_17_ ( .PAD(pad[17]), .C(in[17]), .OEN(oen[17]),
     .I(out[17]), .REN(ren[17]));
PDUW08DGZ I98_16_ ( .PAD(pad[16]), .C(in[16]), .OEN(oen[16]),
     .I(out[16]), .REN(ren[16]));
PDUW08DGZ I98_15_ ( .PAD(pad[15]), .C(in[15]), .OEN(oen[15]),
     .I(out[15]), .REN(ren[15]));
PDUW08DGZ I65_9_ ( .PAD(pad[9]), .C(in[9]), .OEN(oen[9]), .I(out[9]),
     .REN(ren[9]));
PDUW08DGZ I65_8_ ( .PAD(pad[8]), .C(in[8]), .OEN(oen[8]), .I(out[8]),
     .REN(ren[8]));
PDUW08DGZ I62_14_ ( .PAD(pad[14]), .C(in[14]), .OEN(oen[14]),
     .I(out[14]), .REN(ren[14]));
PDUW08DGZ I62_13_ ( .PAD(pad[13]), .C(in[13]), .OEN(oen[13]),
     .I(out[13]), .REN(ren[13]));
PDUW08DGZ I62_12_ ( .PAD(pad[12]), .C(in[12]), .OEN(oen[12]),
     .I(out[12]), .REN(ren[12]));
PDUW08DGZ I62_11_ ( .PAD(pad[11]), .C(in[11]), .OEN(oen[11]),
     .I(out[11]), .REN(ren[11]));
PDUW08DGZ I62_10_ ( .PAD(pad[10]), .C(in[10]), .OEN(oen[10]),
     .I(out[10]), .REN(ren[10]));
PDT08DGZ I42 ( .OEN(tdo_en), .I(tdo_int), .PAD(Tdo));
PDIDGZ I55 ( .PAD(Tdi), .C(tdi_int));
PDIDGZ I40 ( .C(tck_int), .PAD(Tck));
PDIDGZ I41 ( .C(trstb_int), .PAD(TRSTb));
PDIDGZ I39 ( .C(tms_int), .PAD(Tms));
PVSS3DGZ I85_1_ ( .VSS(gnd_));
PVSS3DGZ I85_0_ ( .VSS(gnd_));
PVSS3DGZ I93_2_ ( .VSS(gnd_));
PVSS3DGZ I93_1_ ( .VSS(gnd_));
PVSS3DGZ I93_0_ ( .VSS(gnd_));
PVSS3DGZ I97_1_ ( .VSS(gnd_));
PVSS3DGZ I97_0_ ( .VSS(gnd_));
PVSS3DGZ I96_1_ ( .VSS(gnd_));
PVSS3DGZ I96_0_ ( .VSS(gnd_));
PVDD1DGZ I72_1_ ( .VDD(vdd_));
PVDD1DGZ I72_0_ ( .VDD(vdd_));
PVDD2POC I82 ( .VDDPST(vddp_));
PVDD2POC I79 ( .VDDPST(vddio_rightbank));
PVDD2DGZ I91_1_ ( .VDDPST(vddio_rightbank));
PVDD2DGZ I91_0_ ( .VDDPST(vddio_rightbank));
PVDD2DGZ I78 ( .VDDPST(vddio_rightbank));
PVDD2DGZ I95_1_ ( .VDDPST(vddio_rightbank));
PVDD2DGZ I95_0_ ( .VDDPST(vddio_rightbank));

endmodule
// Library - NVCM, Cell - ml_core_ctrl_top, View - schematic
// LAST TIME SAVED: May  4 14:26:28 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_ctrl_top ( gwl_b_gnden_25, nv_dataout, yp1, yp1_b_25,
     yp2, yp2_b_25, yp3_25, yp3_b_25, yp_test, yp_test_25,
     yp_test_b_25, bl_out, bl_pgm_glb, s_b_25, s_b_hv, sb25sup_25,
     sbhvsup_hv, vblinhi_pgm_25, vdd_tieh, vpxa, ysup_25, dec_ok_25,
     fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, tm_allbl_h, tm_allbl_l, tm_allwl_h,
     tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr );
output  gwl_b_gnden_25, nv_dataout;

inout  bl_out, bl_pgm_glb, sb25sup_25, sbhvsup_hv, vblinhi_pgm_25,
     vdd_tieh, vpxa, ysup_25;

input  dec_ok_25, fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, saen_25, saen_b_vpxa, testdec_en_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [1:0]  yp_test_b_25;
output [1:0]  yp_test;
output [1:0]  yp_test_25;
output [5:0]  yp1_b_25;
output [7:0]  yp3_25;
output [5:0]  yp1;
output [7:0]  yp2_b_25;
output [7:0]  yp3_b_25;
output [7:0]  yp2;

inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefpgm;
input [4:1]  sa_pgate_vpxa;
input [4:1]  sa_ngate_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  sb25_gnd_25;

wire  [3:0]  sbhv_gnd_25;

wire  [3:0]  sbhv_high_25;

wire  [3:0]  sb25_high_25;

wire  [7:5]  dec_trim;

wire  [7:0]  yp3_sel;

wire  [7:0]  yp2_sel;

wire  [5:0]  yp1_sel;



inv_25 I38 ( .IN(net293), .OUT(gwl_b_gnden_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I30 ( .IN(fsm_gwlbdis_b_25), .OUT(net293), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_core_ctrl_logic Icore_ctrl_logic ( .yp1_sel(yp1_sel[5:0]),
     .yp2_sel(yp2_sel[7:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_tm_allwl_l(tm_allwl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25), .tm_tcol(tm_tcol),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_allbl_l(tm_allbl_l), .fsm_pgm(fsm_pgm),
     .fsm_tm_allbl_h(tm_allbl_h), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_nvcmen(fsm_nvcmen), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd(fsm_blkadd[3:0]), .yp_test(yp_test[1:0]),
     .yp21_b_low_b(yp21_b_low_b), .yp3_sel(yp3_sel[7:0]),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .sbhv_high_25(sbhv_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sb25_gnd_25(sb25_gnd_25[3:0]),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .dec_trim(dec_trim[7:5]));
vdd_tiehigh I117_9_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_8_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_7_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_6_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_5_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_4_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_3_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_2_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_1_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_0_ ( .vdd_tieh(vdd_tieh));
ml_core_sa_top Icore_sa_top ( .tm_dma(tm_dma),
     .fsm_tm_testdec(fsm_tm_testdec), .tm_testdec_wr(tm_testdec_wr),
     .testdec_en_b_25(testdec_en_b_25), .dec_ok_25(dec_ok_25),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .dec_trim(dec_trim[7:5]),
     .nv_dataout(nv_dataout), .vpxa(vpxa), .bl_pgm_glb(bl_pgm_glb),
     .bl_out(bl_out));
ml_wp_ctrl Iml_wp_ctrl ( .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .sbhv_high_25(sbhv_high_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_gnd_25(sb25_gnd_25[3:0]), .s_b_25(s_b_25[3:0]),
     .s_b_hv(s_b_hv[3:0]));
ml_ymux_ctrl Iml_ymux_ctrl ( .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]),
     .yp1(yp1[5:0]), .yp1_b_25(yp1_b_25[5:0]), .yp2_sel(yp2_sel[7:0]),
     .yp1_sel(yp1_sel[5:0]), .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_sel(yp3_sel[7:0]), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test_b_high_b(gnd_),
     .yp_test_b_low_b(gnd_), .yp_test(yp_test[1:0]),
     .yp2_b_low_b(yp21_b_low_b), .yp1_b_low_b(yp21_b_low_b),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .yp_test_25(yp_test_25[1:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_testdec_bgen, View - schematic
// LAST TIME SAVED: Jan 21 10:19:00 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_testdec_bgen ( dec_ok_25, dec_bias_25, dec_det_25,
     testdec_en_b_25, testdec_prec_b_25 );
output  dec_ok_25;

inout  dec_bias_25, dec_det_25;

input  testdec_en_b_25, testdec_prec_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I38 ( .IN(dec_det_25), .OUT(dec_ok_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M23 ( .D(dec_det_25), .B(vddp_), .G(testdec_prec_b_25),
     .S(vddp_));
pch_25  M18_1_ ( .D(dec_bias_sup), .B(vddp_), .G(testdec_en_b_25),
     .S(vddp_));
pch_25  M18_0_ ( .D(dec_bias_sup), .B(vddp_), .G(testdec_en_b_25),
     .S(vddp_));
pch_25  M16 ( .D(net049), .B(vddp_), .G(testdec_en_b_25), .S(vddp_));
pch_25  M19 ( .D(ngate), .B(vddp_), .G(dec_bias_25), .S(net049));
pch_25  M8 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
pch_25  M9_1_ ( .D(dec_det_25), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
pch_25  M9_0_ ( .D(dec_det_25), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
nch_25  M14 ( .D(ngate), .B(GND_), .G(dec_bias_25), .S(gnd_));
nch_25  M15 ( .D(ngate), .B(GND_), .G(testdec_en_b_25), .S(gnd_));
nch_25  M10 ( .D(dec_bias_sup), .B(GND_), .G(ngate), .S(dec_bias_25));
nch_25  M13 ( .D(dec_bias_25), .B(GND_), .G(testdec_en_b_25),
     .S(gnd_));
nch_25  M4 ( .D(dec_det_25), .B(GND_), .G(testdec_en_b_25), .S(gnd_));
nch_25  M17 ( .D(dec_bias_25), .B(GND_), .G(dec_bias_25), .S(gnd_));
nch_25  M20 ( .D(dec_bias_p), .B(GND_), .G(dec_bias_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_testdec_columns, View - schematic
// LAST TIME SAVED: Feb 26 14:35:47 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_testdec_columns ( bl, dec_det_even_25, dec_det_odd_25 );

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(vdd_), .B(gnd_), .G(dec_det_even_25), .S(bl[0]));
nch_25  M4 ( .D(vdd_), .B(gnd_), .G(dec_det_odd_25), .S(bl[1]));

endmodule
// Library - NVCM, Cell - ml_testdec_columnsx330, View - schematic
// LAST TIME SAVED: Feb 26 14:35:34 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_testdec_columnsx330 ( bl, bl_dummyl, bl_dummyr, bl_test,
     dec_det_even_25, dec_det_odd_25 );

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl_dummyl;
inout [327:0]  bl;
inout [1:0]  bl_dummyr;
inout [1:0]  bl_test;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_testdec_columns Itestdec_columns_dml (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyl[1:0]));
ml_testdec_columns Itestdec_columns_163_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[327:326]));
ml_testdec_columns Itestdec_columns_162_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[325:324]));
ml_testdec_columns Itestdec_columns_161_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[323:322]));
ml_testdec_columns Itestdec_columns_160_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[321:320]));
ml_testdec_columns Itestdec_columns_159_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[319:318]));
ml_testdec_columns Itestdec_columns_158_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[317:316]));
ml_testdec_columns Itestdec_columns_157_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[315:314]));
ml_testdec_columns Itestdec_columns_156_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[313:312]));
ml_testdec_columns Itestdec_columns_155_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[311:310]));
ml_testdec_columns Itestdec_columns_154_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[309:308]));
ml_testdec_columns Itestdec_columns_153_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[307:306]));
ml_testdec_columns Itestdec_columns_152_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[305:304]));
ml_testdec_columns Itestdec_columns_151_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[303:302]));
ml_testdec_columns Itestdec_columns_150_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[301:300]));
ml_testdec_columns Itestdec_columns_149_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[299:298]));
ml_testdec_columns Itestdec_columns_148_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[297:296]));
ml_testdec_columns Itestdec_columns_147_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[295:294]));
ml_testdec_columns Itestdec_columns_146_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[293:292]));
ml_testdec_columns Itestdec_columns_145_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[291:290]));
ml_testdec_columns Itestdec_columns_144_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[289:288]));
ml_testdec_columns Itestdec_columns_143_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[287:286]));
ml_testdec_columns Itestdec_columns_142_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[285:284]));
ml_testdec_columns Itestdec_columns_141_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[283:282]));
ml_testdec_columns Itestdec_columns_140_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[281:280]));
ml_testdec_columns Itestdec_columns_139_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[279:278]));
ml_testdec_columns Itestdec_columns_138_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[277:276]));
ml_testdec_columns Itestdec_columns_137_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[275:274]));
ml_testdec_columns Itestdec_columns_136_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[273:272]));
ml_testdec_columns Itestdec_columns_135_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[271:270]));
ml_testdec_columns Itestdec_columns_134_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[269:268]));
ml_testdec_columns Itestdec_columns_133_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[267:266]));
ml_testdec_columns Itestdec_columns_132_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[265:264]));
ml_testdec_columns Itestdec_columns_131_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[263:262]));
ml_testdec_columns Itestdec_columns_130_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[261:260]));
ml_testdec_columns Itestdec_columns_129_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[259:258]));
ml_testdec_columns Itestdec_columns_128_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[257:256]));
ml_testdec_columns Itestdec_columns_127_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[255:254]));
ml_testdec_columns Itestdec_columns_126_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[253:252]));
ml_testdec_columns Itestdec_columns_125_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[251:250]));
ml_testdec_columns Itestdec_columns_124_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[249:248]));
ml_testdec_columns Itestdec_columns_123_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[247:246]));
ml_testdec_columns Itestdec_columns_122_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[245:244]));
ml_testdec_columns Itestdec_columns_121_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[243:242]));
ml_testdec_columns Itestdec_columns_120_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[241:240]));
ml_testdec_columns Itestdec_columns_119_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[239:238]));
ml_testdec_columns Itestdec_columns_118_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[237:236]));
ml_testdec_columns Itestdec_columns_117_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[235:234]));
ml_testdec_columns Itestdec_columns_116_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[233:232]));
ml_testdec_columns Itestdec_columns_115_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[231:230]));
ml_testdec_columns Itestdec_columns_114_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[229:228]));
ml_testdec_columns Itestdec_columns_113_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[227:226]));
ml_testdec_columns Itestdec_columns_112_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[225:224]));
ml_testdec_columns Itestdec_columns_111_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[223:222]));
ml_testdec_columns Itestdec_columns_110_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[221:220]));
ml_testdec_columns Itestdec_columns_109_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[219:218]));
ml_testdec_columns Itestdec_columns_108_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[217:216]));
ml_testdec_columns Itestdec_columns_107_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[215:214]));
ml_testdec_columns Itestdec_columns_106_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[213:212]));
ml_testdec_columns Itestdec_columns_105_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[211:210]));
ml_testdec_columns Itestdec_columns_104_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[209:208]));
ml_testdec_columns Itestdec_columns_103_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[207:206]));
ml_testdec_columns Itestdec_columns_102_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[205:204]));
ml_testdec_columns Itestdec_columns_101_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[203:202]));
ml_testdec_columns Itestdec_columns_100_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[201:200]));
ml_testdec_columns Itestdec_columns_99_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[199:198]));
ml_testdec_columns Itestdec_columns_98_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[197:196]));
ml_testdec_columns Itestdec_columns_97_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[195:194]));
ml_testdec_columns Itestdec_columns_96_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[193:192]));
ml_testdec_columns Itestdec_columns_95_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[191:190]));
ml_testdec_columns Itestdec_columns_94_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[189:188]));
ml_testdec_columns Itestdec_columns_93_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[187:186]));
ml_testdec_columns Itestdec_columns_92_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[185:184]));
ml_testdec_columns Itestdec_columns_91_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[183:182]));
ml_testdec_columns Itestdec_columns_90_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[181:180]));
ml_testdec_columns Itestdec_columns_89_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[179:178]));
ml_testdec_columns Itestdec_columns_88_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[177:176]));
ml_testdec_columns Itestdec_columns_87_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[175:174]));
ml_testdec_columns Itestdec_columns_86_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[173:172]));
ml_testdec_columns Itestdec_columns_85_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[171:170]));
ml_testdec_columns Itestdec_columns_84_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[169:168]));
ml_testdec_columns Itestdec_columns_83_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[167:166]));
ml_testdec_columns Itestdec_columns_82_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[165:164]));
ml_testdec_columns Itestdec_columns_81_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[163:162]));
ml_testdec_columns Itestdec_columns_80_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[161:160]));
ml_testdec_columns Itestdec_columns_79_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[159:158]));
ml_testdec_columns Itestdec_columns_78_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[157:156]));
ml_testdec_columns Itestdec_columns_77_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[155:154]));
ml_testdec_columns Itestdec_columns_76_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[153:152]));
ml_testdec_columns Itestdec_columns_75_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[151:150]));
ml_testdec_columns Itestdec_columns_74_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[149:148]));
ml_testdec_columns Itestdec_columns_73_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[147:146]));
ml_testdec_columns Itestdec_columns_72_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[145:144]));
ml_testdec_columns Itestdec_columns_71_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[143:142]));
ml_testdec_columns Itestdec_columns_70_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[141:140]));
ml_testdec_columns Itestdec_columns_69_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[139:138]));
ml_testdec_columns Itestdec_columns_68_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[137:136]));
ml_testdec_columns Itestdec_columns_67_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[135:134]));
ml_testdec_columns Itestdec_columns_66_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[133:132]));
ml_testdec_columns Itestdec_columns_65_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[131:130]));
ml_testdec_columns Itestdec_columns_64_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[129:128]));
ml_testdec_columns Itestdec_columns_63_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[127:126]));
ml_testdec_columns Itestdec_columns_62_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[125:124]));
ml_testdec_columns Itestdec_columns_61_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[123:122]));
ml_testdec_columns Itestdec_columns_60_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[121:120]));
ml_testdec_columns Itestdec_columns_59_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[119:118]));
ml_testdec_columns Itestdec_columns_58_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[117:116]));
ml_testdec_columns Itestdec_columns_57_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[115:114]));
ml_testdec_columns Itestdec_columns_56_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[113:112]));
ml_testdec_columns Itestdec_columns_55_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[111:110]));
ml_testdec_columns Itestdec_columns_54_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[109:108]));
ml_testdec_columns Itestdec_columns_53_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[107:106]));
ml_testdec_columns Itestdec_columns_52_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[105:104]));
ml_testdec_columns Itestdec_columns_51_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[103:102]));
ml_testdec_columns Itestdec_columns_50_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[101:100]));
ml_testdec_columns Itestdec_columns_49_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[99:98]));
ml_testdec_columns Itestdec_columns_48_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[97:96]));
ml_testdec_columns Itestdec_columns_47_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[95:94]));
ml_testdec_columns Itestdec_columns_46_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[93:92]));
ml_testdec_columns Itestdec_columns_45_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[91:90]));
ml_testdec_columns Itestdec_columns_44_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[89:88]));
ml_testdec_columns Itestdec_columns_43_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[87:86]));
ml_testdec_columns Itestdec_columns_42_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[85:84]));
ml_testdec_columns Itestdec_columns_41_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[83:82]));
ml_testdec_columns Itestdec_columns_40_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[81:80]));
ml_testdec_columns Itestdec_columns_39_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[79:78]));
ml_testdec_columns Itestdec_columns_38_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[77:76]));
ml_testdec_columns Itestdec_columns_37_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[75:74]));
ml_testdec_columns Itestdec_columns_36_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[73:72]));
ml_testdec_columns Itestdec_columns_35_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[71:70]));
ml_testdec_columns Itestdec_columns_34_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[69:68]));
ml_testdec_columns Itestdec_columns_33_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[67:66]));
ml_testdec_columns Itestdec_columns_32_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[65:64]));
ml_testdec_columns Itestdec_columns_31_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[63:62]));
ml_testdec_columns Itestdec_columns_30_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[61:60]));
ml_testdec_columns Itestdec_columns_29_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[59:58]));
ml_testdec_columns Itestdec_columns_28_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[57:56]));
ml_testdec_columns Itestdec_columns_27_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[55:54]));
ml_testdec_columns Itestdec_columns_26_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[53:52]));
ml_testdec_columns Itestdec_columns_25_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[51:50]));
ml_testdec_columns Itestdec_columns_24_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[49:48]));
ml_testdec_columns Itestdec_columns_23_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[47:46]));
ml_testdec_columns Itestdec_columns_22_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[45:44]));
ml_testdec_columns Itestdec_columns_21_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[43:42]));
ml_testdec_columns Itestdec_columns_20_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[41:40]));
ml_testdec_columns Itestdec_columns_19_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[39:38]));
ml_testdec_columns Itestdec_columns_18_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[37:36]));
ml_testdec_columns Itestdec_columns_17_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[35:34]));
ml_testdec_columns Itestdec_columns_16_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[33:32]));
ml_testdec_columns Itestdec_columns_15_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[31:30]));
ml_testdec_columns Itestdec_columns_14_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[29:28]));
ml_testdec_columns Itestdec_columns_13_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[27:26]));
ml_testdec_columns Itestdec_columns_12_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[25:24]));
ml_testdec_columns Itestdec_columns_11_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[23:22]));
ml_testdec_columns Itestdec_columns_10_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[21:20]));
ml_testdec_columns Itestdec_columns_9_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[19:18]));
ml_testdec_columns Itestdec_columns_8_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[17:16]));
ml_testdec_columns Itestdec_columns_7_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[15:14]));
ml_testdec_columns Itestdec_columns_6_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[13:12]));
ml_testdec_columns Itestdec_columns_5_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[11:10]));
ml_testdec_columns Itestdec_columns_4_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[9:8]));
ml_testdec_columns Itestdec_columns_3_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[7:6]));
ml_testdec_columns Itestdec_columns_2_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[5:4]));
ml_testdec_columns Itestdec_columns_1_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[3:2]));
ml_testdec_columns Itestdec_columns_0_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[1:0]));
ml_testdec_columns Itestdec_columns_dmr (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyr[1:0]));
ml_testdec_columns Itestdec_columns_tst (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_test[1:0]));

endmodule
// Library - NVCM, Cell - ml_ymux_yp3_x8, View - schematic
// LAST TIME SAVED: Feb 26 14:33:55 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_yp3_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M5_7_ ( .D(bl[7]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_6_ ( .D(bl[6]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_5_ ( .D(bl[5]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_4_ ( .D(bl[4]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_3_ ( .D(bl[3]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_2_ ( .D(bl[2]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_1_ ( .D(bl[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_0_ ( .D(bl[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
nch_25  M22 ( .D(bl[6]), .B(GND_), .G(yp3_25[6]), .S(bl_out));
nch_25  M1 ( .D(bl[4]), .B(GND_), .G(yp3_25[4]), .S(bl_out));
nch_25  M24 ( .D(bl[2]), .B(GND_), .G(yp3_25[2]), .S(bl_out));
nch_25  M25 ( .D(bl[0]), .B(GND_), .G(yp3_25[0]), .S(bl_out));
nch_25  M26 ( .D(bl[0]), .B(GND_), .G(yp3_b_25[0]), .S(vblinhi_rde));
nch_25  M27 ( .D(bl[1]), .B(GND_), .G(yp3_b_25[1]), .S(vblinhi_rdo));
nch_25  M28 ( .D(bl[1]), .B(GND_), .G(yp3_25[1]), .S(bl_out));
nch_25  M29 ( .D(bl[3]), .B(GND_), .G(yp3_b_25[3]), .S(vblinhi_rdo));
nch_25  M30 ( .D(bl[3]), .B(GND_), .G(yp3_25[3]), .S(bl_out));
nch_25  M31 ( .D(bl[2]), .B(GND_), .G(yp3_b_25[2]), .S(vblinhi_rde));
nch_25  M20 ( .D(bl[4]), .B(GND_), .G(yp3_b_25[4]), .S(vblinhi_rde));
nch_25  M19 ( .D(bl[5]), .B(GND_), .G(yp3_b_25[5]), .S(vblinhi_rdo));
nch_25  M21 ( .D(bl[5]), .B(GND_), .G(yp3_25[5]), .S(bl_out));
nch_25  M13 ( .D(bl[7]), .B(GND_), .G(yp3_b_25[7]), .S(vblinhi_rdo));
nch_25  M23 ( .D(bl[7]), .B(GND_), .G(yp3_25[7]), .S(bl_out));
nch_25  M18 ( .D(bl[6]), .B(GND_), .G(yp3_b_25[6]), .S(vblinhi_rde));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x8, View - schematic
// LAST TIME SAVED: May  4 13:03:21 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_bls_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_dummy, View - schematic
// LAST TIME SAVED: Feb 26 14:34:35 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_bls_dummy ( bl_dummyr, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, pgminhi_dmmy_b_25, vdd_tieh );
inout  vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo;

input  pgminhi_dmmy_b_25, vdd_tieh;

inout [1:0]  bl_dummyr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(bl_dummyr[1]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rdo));
nch_25  M18 ( .D(bl_dummyr[0]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rde));
pch_25  M8 ( .D(bl_dummyr[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M0 ( .D(bl_dummyr[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_yp2_8, View - schematic
// LAST TIME SAVED: Feb 12 15:37:16 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_yp2_8 ( bl, bl_out, vblinhi_rde, vblinhi_rdo, yp2,
     yp2_b_25 );
inout  bl_out, vblinhi_rde, vblinhi_rdo;


inout [7:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M17 ( .D(bl[7]), .B(GND_), .G(yp2_b_25[7]), .S(vblinhi_rdo));
nch_25  M16 ( .D(bl[6]), .B(GND_), .G(yp2_b_25[6]), .S(vblinhi_rde));
nch_25  M11 ( .D(bl[1]), .B(GND_), .G(yp2_b_25[1]), .S(vblinhi_rdo));
nch_25  M20 ( .D(bl[0]), .B(GND_), .G(yp2_b_25[0]), .S(vblinhi_rde));
nch_25  M15 ( .D(bl[5]), .B(GND_), .G(yp2_b_25[5]), .S(vblinhi_rdo));
nch_25  M14 ( .D(bl[4]), .B(GND_), .G(yp2_b_25[4]), .S(vblinhi_rde));
nch_25  M13 ( .D(bl[3]), .B(GND_), .G(yp2_b_25[3]), .S(vblinhi_rdo));
nch_25  M12 ( .D(bl[2]), .B(GND_), .G(yp2_b_25[2]), .S(vblinhi_rde));
nch_hvt  M3 ( .D(bl[3]), .B(GND_), .G(yp2[3]), .S(bl_out));
nch_hvt  M1 ( .D(bl[2]), .B(GND_), .G(yp2[2]), .S(bl_out));
nch_hvt  M0 ( .D(bl[1]), .B(GND_), .G(yp2[1]), .S(bl_out));
nch_hvt  M7 ( .D(bl[7]), .B(GND_), .G(yp2[7]), .S(bl_out));
nch_hvt  M6 ( .D(bl[6]), .B(GND_), .G(yp2[6]), .S(bl_out));
nch_hvt  M5 ( .D(bl[5]), .B(GND_), .G(yp2[5]), .S(bl_out));
nch_hvt  M2 ( .D(bl[0]), .B(GND_), .G(yp2[0]), .S(bl_out));
nch_hvt  M4 ( .D(bl[4]), .B(GND_), .G(yp2[4]), .S(bl_out));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x64, View - schematic
// LAST TIME SAVED: Feb 26 14:34:16 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_bls_x64 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp2, yp2_b_25, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [63:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
input [7:0]  yp3_25;
input [7:0]  yp3_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  bl_med;



ml_ymux_yp2_8 Iml_ymux_yp2_x8 ( .bl(bl_med[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[0]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_2 ( .vdd_tieh(vdd_tieh), .bl(bl[23:16]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[2]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_3 ( .vdd_tieh(vdd_tieh), .bl(bl[31:24]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[3]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_6 ( .vdd_tieh(vdd_tieh), .bl(bl[55:48]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[6]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_7 ( .vdd_tieh(vdd_tieh), .bl(bl[63:56]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[7]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_5 ( .vdd_tieh(vdd_tieh), .bl(bl[47:40]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[5]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_4 ( .vdd_tieh(vdd_tieh), .bl(bl[39:32]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[4]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_1 ( .vdd_tieh(vdd_tieh), .bl(bl[15:8]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[1]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x328, View - schematic
// LAST TIME SAVED: May  4 14:26:48 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_bls_x328 ( bl, bl_dummyl, bl_dummyr, bl_out, bl_test,
     vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh,
     pgminhi_dmmy_b_25, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25,
     yp_test, yp_test_25, yp_test_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25;

inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;
inout [1:0]  bl_dummyr;
inout [327:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp2_b_25;
input [7:0]  yp2;
input [1:0]  yp_test_b_25;
input [5:0]  yp1_b_25;
input [1:0]  yp_test_25;
input [7:0]  yp3_25;
input [1:0]  yp_test;
input [5:0]  yp1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:5]  blx8_out;

wire  [0:4]  blx64_out;



ml_ymux_bls_x8 Iml_ymux_bls_x8 ( .bl_out(blx8_out[5]),
     .bl(bl[327:320]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_r ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyr[1:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_l ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyl[1:0]));
pch_25  M7 ( .D(bl_test[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M8 ( .D(bl_test[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
ml_ymux_bls_x64 Iml_ymux_bls_x64_0 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[0]), .bl(bl[63:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_2 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[2]), .bl(bl[191:128]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_4 ( .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]), .bl(bl[319:256]),
     .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]), .bl_out(blx64_out[4]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo));
ml_ymux_bls_x64 Iml_ymux_bls_x64_1 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[1]), .bl(bl[127:64]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_3 ( .yp2(yp2[7:0]), .bl_out(blx64_out[3]),
     .bl(bl[255:192]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .yp2_b_25(yp2_b_25[7:0]), .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]));
nch_hvt  M21 ( .D(net224), .B(GND_), .G(yp_test[1]), .S(bl_out));
nch_hvt  M19 ( .D(net228), .B(GND_), .G(yp_test[1]), .S(net224));
nch_hvt  M23 ( .D(net232), .B(GND_), .G(yp_test[0]), .S(bl_out));
nch_hvt  M28 ( .D(net236), .B(GND_), .G(yp1[5]), .S(bl_out));
nch_hvt  M0 ( .D(blx64_out[2]), .B(GND_), .G(yp1[2]), .S(bl_out));
nch_hvt  M22 ( .D(net244), .B(GND_), .G(yp_test[0]), .S(net232));
nch_hvt  M24 ( .D(blx64_out[0]), .B(GND_), .G(yp1[0]), .S(bl_out));
nch_hvt  M30 ( .D(blx8_out[5]), .B(GND_), .G(yp1[5]), .S(net236));
nch_hvt  M3 ( .D(blx64_out[4]), .B(GND_), .G(yp1[4]), .S(bl_out));
nch_hvt  M4 ( .D(blx64_out[3]), .B(GND_), .G(yp1[3]), .S(bl_out));
nch_hvt  M2 ( .D(blx64_out[1]), .B(GND_), .G(yp1[1]), .S(bl_out));
nch_25  M27 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[0]),
     .S(blx64_out[0]));
nch_25  M26 ( .D(vblinhi_rdo), .B(GND_), .G(yp_test_b_25[1]),
     .S(bl_test[1]));
nch_25  M25 ( .D(bl_test[1]), .B(GND_), .G(yp_test_25[1]), .S(net228));
nch_25  M18 ( .D(vblinhi_rde), .B(GND_), .G(yp_test_b_25[0]),
     .S(bl_test[0]));
nch_25  M29 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[5]),
     .S(blx8_out[5]));
nch_25  M17 ( .D(bl_test[0]), .B(GND_), .G(yp_test_25[0]), .S(net244));
nch_25  M1 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[2]),
     .S(blx64_out[2]));
nch_25  M20 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[1]),
     .S(blx64_out[1]));
nch_25  M5 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[4]),
     .S(blx64_out[4]));
nch_25  M6 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[3]),
     .S(blx64_out[3]));

endmodule
// Library - sbtlibn65lp, Cell - vddp_tiehigh, View - schematic
// LAST TIME SAVED: May  8 16:23:22 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module vddp_tiehigh ( vddp_tieh );
inout  vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M8 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net9), .S(vddp_));

endmodule
// Library - NVCM, Cell - ml_core_338x112_top_1f, View - schematic
// LAST TIME SAVED: Feb  9 11:10:00 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_338x112_top_1f ( nv_dataout, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25,
     sa_ngate_25, sa_pgate_vpxa, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr, wr );
output  nv_dataout;

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     pgminhi_dmmy_b_25, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

input [4:1]  sa_ngate_25;
input [3:0]  fsm_blkadd;
input [26:0]  gwp_hv;
input [107:0]  wr;
input [4:1]  sa_pgate_vpxa;
input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefpgm;
input [26:0]  gwl_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_b_25;

wire  [5:0]  yp1;

wire  [5:0]  yp1_b_25;

wire  [1:0]  bl_dummyr;

wire  [327:0]  bl;

wire  [7:0]  yp2;

wire  [1:0]  yp_test;

wire  [7:0]  yp3_b_25;

wire  [107:0]  wp;

wire  [1:0]  yp_test_b_25;

wire  [7:0]  yp2_b_25;

wire  [1:0]  bl_dummyl;

wire  [1:0]  bl_test;

wire  [3:0]  s_b_hv;

wire  [1:0]  yp_test_25;

wire  [7:0]  yp3;



ml_core_sa_spare Iml_core_sa_spare ( );
ml_testdec_rowsx108_1f Iml_testdec_rowsx108_1f ( .wp(wp[107:0]),
     .wr(wr[107:0]), .dec_bias_25(dec_bias), .dec_det_25(dec_det_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25));
ml_rock_lwldrv_wp_x108_1f Iml_rock_lwldrv_wp_x108_1f ( .wp(wp[107:0]),
     .gwl_b_25(gwl_b_25[26:0]), .gwp_hv(gwp_hv[26:0]),
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .ngate_25(ngate_25));
nvcm_cell_338x112_1f Invcm_cell_338x112_1f ( .wp(wp[107:0]),
     .wr(wr[107:0]), .bl_dummyr(bl_dummyr[1:0]), .wr_dummyt({net156,
     net156}), .wr_dummyb({net156, net156}), .wp_dummyt({net156,
     net156}), .wp_dummyb({net156, net156}), .bl_test(bl_test[1:0]),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
vdd_tielow I47 ( .gnd_tiel(net156));
inv_hvt I131 ( .A(nv_dataout_in), .Y(net158));
inv_hvt I45 ( .A(net158), .Y(nv_dataout));
ml_core_ctrl_top Icore_ctrl_top ( .yp2_b_25(yp2_b_25[7:0]),
     .yp2(yp2[7:0]), .yp1_b_25(yp1_b_25[5:0]), .yp1(yp1[5:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .gwl_b_gnden_25(gwl_b_gnden_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .vdd_tieh(vdd_tieh), .tm_testdec_wr(tm_testdec_wr),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .testdec_en_b_25(testdec_en_b_25),
     .saen_b_vpxa(saen_b_vpxa), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .dec_ok_25(dec_ok_25), .yp_test_b_25(yp_test_b_25[1:0]),
     .yp_test_25(yp_test_25[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .nv_dataout(nv_dataout_in), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_pgm_25(vblinhi_pgm_25),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .bl_out(bl_out),
     .yp_test(yp_test[1:0]));
ml_testdec_bgen Itestdec_bgen ( .dec_ok_25(dec_ok_25),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25), .dec_det_25(dec_det_25),
     .dec_bias_25(dec_bias));
ml_testdec_columnsx330 Itestdec_columnsx330 (
     .bl_dummyr(bl_dummyr[1:0]), .bl_dummyl(bl_dummyl[1:0]),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[327:0]),
     .bl_test(bl_test[1:0]));
ml_ymux_bls_x328 Iml_ymux_bls_x328 ( .yp1_b_25(yp1_b_25[5:0]),
     .yp1(yp1[5:0]), .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]),
     .vdd_tieh(vdd_tieh), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .bl_dummyl(bl_dummyl[1:0]), .bl_dummyr(bl_dummyr[1:0]),
     .bl_test(bl_test[1:0]), .yp_test_b_25(yp_test_b_25[1:0]),
     .yp_test_25(yp_test_25[1:0]), .yp_test(yp_test[1:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3[7:0]),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .vblinhi_pgm_25(vblinhi_pgm_25), .bl_out(bl_out), .bl(bl[327:0]));

endmodule
// Library - NVCM, Cell - ml_core_bank_0_1f, View - schematic
// LAST TIME SAVED: Mar  5 15:01:51 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_bank_0_1f ( nv_dataout, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv,
     pgminhi_dmmy_b_25, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     pgminhi_dmmy_b_25, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [3:0]  nv_dataout;

input [4:1]  sa_pgate_vpxa;
input [2:0]  fsm_trim_rrefpgm;
input [26:0]  gwp_hv;
input [4:1]  sa_ngate_25;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefrd;
input [1:0]  fsm_rowadd;
input [107:0]  wr;
input [3:0]  fsm_blkadd;
input [3:0]  fsm_blkadd_b;
input [26:0]  gwl_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_core_338x112_top_1f blk3 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen), .tm_dma(tm_dma),
     .fsm_tm_trow(fsm_tm_trow), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd[1],
     fsm_blkadd[0]}), .nv_dataout(nv_dataout[3]), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));
ml_core_338x112_top_1f blk1 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen), .tm_dma(tm_dma),
     .fsm_tm_trow(fsm_tm_trow), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd[0]}), .nv_dataout(nv_dataout[1]), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));
ml_core_338x112_top_1f blk2 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen), .tm_dma(tm_dma),
     .fsm_tm_trow(fsm_tm_trow), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd[1],
     fsm_blkadd_b[0]}), .nv_dataout(nv_dataout[2]), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));
ml_core_338x112_top_1f blk0 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen), .tm_dma(tm_dma),
     .fsm_tm_trow(fsm_tm_trow), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd_b[0]}), .nv_dataout(nv_dataout[0]), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));

endmodule
// Library - NVCM, Cell - ml_core_bank_1_1f, View - schematic
// LAST TIME SAVED: Jan 20 11:29:00 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_bank_1_1f ( nv_dataout, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv,
     pgminhi_dmmy_b_25, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     pgminhi_dmmy_b_25, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [8:4]  nv_dataout;

input [107:0]  wr;
input [26:0]  gwp_hv;
input [3:0]  fsm_blkadd;
input [3:0]  fsm_blkadd_b;
input [2:0]  fsm_trim_rrefrd;
input [26:0]  gwl_b_25;
input [8:0]  fsm_coladd;
input [4:1]  sa_ngate_25;
input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefpgm;
input [4:1]  sa_pgate_vpxa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_core_338x112_top_1f blk4 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .nv_dataout(nv_dataout[4]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));
ml_core_338x112_top_1f blk5 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd[0]}),
     .nv_dataout(nv_dataout[5]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));
ml_core_338x112_top_1f blk7 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd[1], fsm_blkadd[0]}),
     .nv_dataout(nv_dataout[7]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));
ml_core_338x112_top_1f blk6 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd[1], fsm_blkadd_b[0]}),
     .nv_dataout(nv_dataout[6]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));
ml_core_338x112_top_1f blk8 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd[3],
     fsm_blkadd_b[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .nv_dataout(nv_dataout[8]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));

endmodule
// Library - NVCM, Cell - ml_core_1f, View - schematic
// LAST TIME SAVED: Jan 20 17:30:10 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_core_1f ( nv_dataout, bgr, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpp_int, vpxa, ysup_25, fsm_blkadd,
     fsm_blkadd_b, fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven,
     fsm_multibl_read, fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_trim_ipp,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo,
     vpp_int, vpxa, ysup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbl_h, tm_allbl_l, tm_allwl_h,
     tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [8:0]  nv_dataout;

input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_trim_rrefpgm;
input [2:0]  fsm_trim_rrefrd;
input [8:0]  fsm_coladd;
input [7:0]  fsm_rowadd;
input [3:0]  fsm_blkadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:1]  sa_ngate_25;

wire  [4:1]  sa_pgate_vpxa;

wire  [26:0]  gwp_hv;

wire  [107:0]  wr;

wire  [26:0]  gwl_b_25;



ml_gwlwr_top_1f Igwlwr_top_1f ( .gwl_b_25(gwl_b_25[26:0]),
     .gwp_hv(gwp_hv[26:0]), .wr(wr[107:0]), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_din(fsm_din), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_wren(fsm_wren), .tm_testdec(fsm_tm_testdec),
     .fsm_tm_allbl_h(tm_allbl_h), .fsm_tm_allwl_l(tm_allwl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .fsm_tm_allbl_l(tm_allbl_l),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_wpen(fsm_wpen),
     .tm_dma(tm_dma), .gwl_b_sup_25(gwl_b_sup_25),
     .tm_testdec_wr(tm_testdec_wr), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wgnden(fsm_wgnden), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .vpxa(vpxa),
     .vpp_int(vpp_int), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr));
ml_core_bank_0_1f bank0_1f ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .ysup_25(ysup_25),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .nv_dataout(nv_dataout[3:0]), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .tm_testdec_wr(tm_testdec_wr));
ml_core_bank_1_1f bank1_1f ( .gwl_b_25(gwl_b_25[26:0]),
     .gwp_hv(gwp_hv[26:0]), .wr(wr[107:0]), .fsm_tm_trow(fsm_tm_trow),
     .tm_dma(tm_dma), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .gwl_b_sup_25(gwl_b_sup_25),
     .ngate_25(ngate_25), .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vpxa(vpxa), .ysup_25(ysup_25),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rst_b(fsm_rst_b),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_wpen(fsm_wpen), .fsm_ymuxdis(fsm_ymuxdis),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]), .saen_25(saen_25),
     .saen_b_vpxa(saen_b_vpxa), .testdec_en_b_25(testdec_en_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_prec_b_25(testdec_prec_b_25), .tm_allbl_h(tm_allbl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd(fsm_blkadd[3:0]),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .nv_dataout(nv_dataout[8:4]),
     .bl_pgm_glb(bl_pgm_glb));

endmodule
// Library - NVCM, Cell - ml_chip_buf, View - schematic
// LAST TIME SAVED: Feb 26 16:35:06 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_chip_buf ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(in), .Y(net120));
inv_hvt I45 ( .A(net120), .Y(out));

endmodule
// Library - NVCM, Cell - ml_chip_buf_top, View - schematic
// LAST TIME SAVED: Apr 21 14:59:16 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_chip_buf_top ( fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_trim_vbg_buf, fsm_vpgmwl_buf,
     fsm_wgnden_buf, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmvfy, fsm_trim_vbg, fsm_vpgmwl, fsm_wgnden );
output  fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf,
     fsm_pgmvfy_buf, fsm_wgnden_buf;

input  fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmvfy,
     fsm_wgnden;

output [2:0]  fsm_vpgmwl_buf;
output [3:0]  fsm_trim_vbg_buf;

input [3:0]  fsm_trim_vbg;
input [2:0]  fsm_vpgmwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_chip_buf I50_2_ ( .in(fsm_vpgmwl[2]), .out(fsm_vpgmwl_buf[2]));
ml_chip_buf I50_1_ ( .in(fsm_vpgmwl[1]), .out(fsm_vpgmwl_buf[1]));
ml_chip_buf I50_0_ ( .in(fsm_vpgmwl[0]), .out(fsm_vpgmwl_buf[0]));
ml_chip_buf I56 ( .in(fsm_wgnden), .out(fsm_wgnden_buf));
ml_chip_buf I49_3_ ( .in(fsm_trim_vbg[3]), .out(fsm_trim_vbg_buf[3]));
ml_chip_buf I49_2_ ( .in(fsm_trim_vbg[2]), .out(fsm_trim_vbg_buf[2]));
ml_chip_buf I49_1_ ( .in(fsm_trim_vbg[1]), .out(fsm_trim_vbg_buf[1]));
ml_chip_buf I49_0_ ( .in(fsm_trim_vbg[0]), .out(fsm_trim_vbg_buf[0]));
ml_chip_buf I51 ( .in(fsm_lshven), .out(fsm_lshven_buf));
ml_chip_buf I53 ( .in(fsm_nvcmen), .out(fsm_nvcmen_buf));
ml_chip_buf I54 ( .in(fsm_pgmdisc), .out(fsm_pgmdisc_buf));
ml_chip_buf I57 ( .in(fsm_pgmvfy), .out(fsm_pgmvfy_buf));
ml_chip_buf I55 ( .in(fsm_pgm), .out(fsm_pgm_buf));

endmodule
// Library - NVCM, Cell - ml_hv2vddp_sw, View - schematic
// LAST TIME SAVED: May  1 11:01:33 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_hv2vddp_sw ( out_hv, hv2vddp, vddp_tieh );
inout  out_hv;

input  hv2vddp, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(sw_vddp_b),
     .sel_25(net035), .out_b_hv(sw_vpp_b), .in_hv(out_hv),
     .vddp_tieh(vddp_tieh));
pch_25  M1 ( .D(net27), .B(out_hv), .G(sw_vpp_b), .S(out_hv));
pch_25  M0 ( .D(net27), .B(vddp_), .G(sw_vddp_b), .S(vddp_));
inv_25 I62 ( .IN(net37), .OUT(sw_vddp_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I71 ( .IN(net060), .OUT(net035), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net060),
     .out_vddio(net37), .in_b(net46));
inv_hvt I65 ( .A(hv2vddp), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));

endmodule
// Library - NVCM, Cell - ml_vpp_ref_sw, View - schematic
// LAST TIME SAVED: Mar 21 16:41:35 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpp_ref_sw ( in, out, sel_b_25 );
inout  in, out;

input  sel_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I281 ( .IN(sel_b_25), .OUT(net122), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nch_25  M12 ( .D(out), .B(GND_), .G(net122), .S(in));
pch_25  M14 ( .D(in), .B(vddp_), .G(sel_b_25), .S(out));

endmodule
// Library - NVCM, Cell - ml_vpp_ref, View - schematic
// LAST TIME SAVED: Apr  7 18:49:59 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpp_ref ( vref_25, bgr, pumpen_25, vppwl_25 );
inout  vref_25;

input  bgr, pumpen_25;

input [2:0]  vppwl_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_b_25;

wire  [7:0]  red_dec_25;



nch_na25  M0 ( .D(net179), .B(GND_), .G(ctrl_gate_25),
     .S(bgr_mirror_25));
nand3_25 I44_7_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[7]),
     .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_6_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[6]),
     .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_5_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[5]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_4_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[4]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_3_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[3]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_2_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[2]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_1_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[1]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_0_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[0]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
ml_vpp_ref_sw I281 ( .in(net92), .out(vref_25),
     .sel_b_25(red_dec_25[6]));
ml_vpp_ref_sw I287 ( .in(net95), .out(vref_25),
     .sel_b_25(red_dec_25[4]));
ml_vpp_ref_sw I283 ( .in(net98), .out(vref_25),
     .sel_b_25(red_dec_25[7]));
ml_vpp_ref_sw I290 ( .in(net0100), .out(vref_25),
     .sel_b_25(red_dec_25[0]));
ml_vpp_ref_sw I288 ( .in(net104), .out(vref_25),
     .sel_b_25(red_dec_25[3]));
ml_vpp_ref_sw I284 ( .in(net139), .out(vref_25),
     .sel_b_25(red_dec_25[5]));
ml_vpp_ref_sw I291 ( .in(net110), .out(vref_25),
     .sel_b_25(red_dec_25[1]));
ml_vpp_ref_sw I292 ( .in(net113), .out(vref_25),
     .sel_b_25(red_dec_25[2]));
// nmoscap_25  C3 ( .MINUS(net0129), .PLUS(net0113));
// nmoscap_25  C2 ( .MINUS(gnd_), .PLUS(ctrl_gate_25));
inv_25 I38 ( .IN(pumpen_25), .OUT(vppref_en_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_2_ ( .IN(vppwl_25[2]), .OUT(vppwl_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_1_ ( .IN(vppwl_25[1]), .OUT(vppwl_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_0_ ( .IN(vppwl_25[0]), .OUT(vppwl_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
rppolywo_m  R11 ( .MINUS(net110), .PLUS(net113), .BULK(GND_));
rppolywo_m  R13 ( .MINUS(net113), .PLUS(net104), .BULK(GND_));
rppolywo_m  R14 ( .MINUS(net113), .PLUS(net104), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(net110), .PLUS(net113), .BULK(GND_));
rppolywo_m  R15 ( .MINUS(net104), .PLUS(net95), .BULK(GND_));
rppolywo_m  R16 ( .MINUS(net104), .PLUS(net95), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net95), .PLUS(net139), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net95), .PLUS(net139), .BULK(GND_));
rppolywo_m  R19 ( .MINUS(net139), .PLUS(net92), .BULK(GND_));
rppolywo_m  R20 ( .MINUS(net139), .PLUS(net92), .BULK(GND_));
rppolywo_m  R21 ( .MINUS(net92), .PLUS(net98), .BULK(GND_));
rppolywo_m  R22 ( .MINUS(net92), .PLUS(net98), .BULK(GND_));
rppolywo_m  R25 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R24 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(net0100), .BULK(GND_));
rppolywo_m  R5 ( .MINUS(net0100), .PLUS(net110), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net0100), .PLUS(net110), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(bgr_mirror_25), .PLUS(net0129), .BULK(GND_));
nch_25  M10 ( .D(net163), .B(GND_), .G(bgr), .S(gnd_));
nch_25  M14 ( .D(net0113), .B(GND_), .G(vppref_en_b_25), .S(gnd_));
nch_25  M15 ( .D(ctrl_gate_25), .B(GND_), .G(vppref_en_b_25),
     .S(gnd_));
nch_25  M8 ( .D(ctrl_gate_25), .B(GND_), .G(bgr_mirror_25),
     .S(net163));
nch_25  M13 ( .D(net0113), .B(GND_), .G(bgr), .S(net163));
pch_25  M18 ( .D(net179), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
pch_25  M5 ( .D(ctrl_gate_25), .B(vddp_), .G(net0113), .S(net175));
pch_25  M6 ( .D(net0113), .B(vddp_), .G(net0113), .S(net175));
pch_25  M7 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));

endmodule
// Library - NVCM, Cell - ml_vpp_ctrl, View - schematic
// LAST TIME SAVED: Apr 30 14:24:32 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpp_ctrl ( pumpen_25, vpint_en, vpp_2_vdd, vppdisc_25,
     vppwl_25, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_vpgmwl_buf, fsm_wgnden );
output  pumpen_25, vpint_en, vpp_2_vdd, vppdisc_25;

input  fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf,
     fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint, fsm_wgnden;

output [2:0]  vppwl_25;

input [2:0]  fsm_vpgmwl_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:2]  net068;

wire  [0:2]  net038;

wire  [0:2]  net082;

wire  [0:2]  net092;



nand4_hvt I75 ( .D(fsm_pgm_buf), .C(fsm_lshven_buf), .A(net0127),
     .Y(net046), .B(net0127));
// nmoscap_25  C7 ( .MINUS(GND_), .PLUS(net0122));
nor2_hvt I111 ( .A(vpp_pumpen_b), .B(net080), .Y(net0133));
nor2_hvt I87 ( .A(vpp_pumpen), .Y(net036), .B(fsm_pgmdisc_buf));
sbtlibn65lp_ml_dff_schematic I77 ( .CLK(net084), .QN(vpp_pumpen_b),
     .R(pgm_dis), .D(vdd_tieh), .Q(vpp_pumpen));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
nand3_hvt I79 ( .C(net086), .A(fsm_pgm_buf), .Y(pgm_dis),
     .B(fsm_nvcmen_buf));
nand2_hvt I104 ( .A(fsm_tm_xforce), .Y(net049), .B(fsm_tm_xvppint));
inv_25 I95_2_ ( .IN(net068[0]), .OUT(vppwl_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_1_ ( .IN(net068[1]), .OUT(vppwl_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_0_ ( .IN(net068[2]), .OUT(vppwl_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I81 ( .IN(net073), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(net088), .OUT(vppdisc_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I96_2_ ( .in(net082[0]), .sup(vddp_),
     .out_vddio_b(net068[0]), .out_vddio(net038[0]), .in_b(net092[0]));
ml_ls_vdd2vdd25 I96_1_ ( .in(net082[1]), .sup(vddp_),
     .out_vddio_b(net068[1]), .out_vddio(net038[1]), .in_b(net092[1]));
ml_ls_vdd2vdd25 I96_0_ ( .in(net082[2]), .sup(vddp_),
     .out_vddio_b(net068[2]), .out_vddio(net038[2]), .in_b(net092[2]));
ml_ls_vdd2vdd25 I84 ( .in(net0133), .sup(vddp_), .out_vddio_b(net073),
     .out_vddio(net074), .in_b(net0134));
ml_ls_vdd2vdd25 I173 ( .in(fsm_pgmdisc_buf), .sup(vddp_),
     .out_vddio_b(net088), .out_vddio(net048), .in_b(net0106));
inv_hvt I107 ( .A(net0122), .Y(net0124));
inv_hvt I109 ( .A(fsm_pgmvfy_buf), .Y(net0127));
inv_hvt I131 ( .A(net049), .Y(net080));
inv_hvt I110_2_ ( .A(net092[0]), .Y(net082[0]));
inv_hvt I110_1_ ( .A(net092[1]), .Y(net082[1]));
inv_hvt I110_0_ ( .A(net092[2]), .Y(net082[2]));
inv_hvt I76 ( .A(net046), .Y(net084));
inv_hvt I108 ( .A(fsm_pgmdisc_buf), .Y(net0122));
inv_hvt I78 ( .A(net0124), .Y(net086));
inv_hvt I113 ( .A(vpp_pumpen_b), .Y(vpint_en));
inv_hvt I91 ( .A(net036), .Y(net089));
inv_hvt I90 ( .A(net089), .Y(vpp_2_vdd));
inv_hvt I98_2_ ( .A(fsm_vpgmwl_buf[2]), .Y(net092[0]));
inv_hvt I98_1_ ( .A(fsm_vpgmwl_buf[1]), .Y(net092[1]));
inv_hvt I98_0_ ( .A(fsm_vpgmwl_buf[0]), .Y(net092[2]));
inv_hvt I112 ( .A(net0133), .Y(net0134));
inv_hvt I101 ( .A(fsm_pgmdisc_buf), .Y(net0106));

endmodule
// Library - misc, Cell - vpp_clamp_finger, View - schematic
// LAST TIME SAVED: Jul 30 12:32:02 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module vpp_clamp_finger ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .B(VSS), .D(net12), .G(VSS), .S(VSS));
nch_25  m1 ( .B(VSS), .D(VPP), .G(VDDIO), .S(net12));

endmodule
// Library - NVCM, Cell - ml_vpp_reg, View - schematic
// LAST TIME SAVED: May  3 15:48:51 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpp_reg ( slow_25, bgr, pbias_25, pump_in, vpp_int,
     pumpen_25, vppdisc_25, vref_25 );
output  slow_25;

inout  bgr, pbias_25, pump_in, vpp_int;

input  pumpen_25, vppdisc_25, vref_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I261 ( .vddp_tieh(net0208));
nch_na25  M11 ( .D(net0199), .B(GND_), .G(vppdisc_25), .S(VDD_));
nch_na25  M22 ( .D(vpp_int), .B(GND_), .G(pump_gate), .S(pump_in));
nch_na25  M1 ( .D(GND_), .B(GND_), .G(pump_gate), .S(GND_));
nch_na25  M10 ( .D(net0203), .B(GND_), .G(net0208), .S(net0199));
nch_na25  M5 ( .D(pump_opamp_out), .B(GND_), .G(vpp_int),
     .S(pump_opamp_out));
inv_25 I211 ( .IN(en_buf_b_25), .OUT(en_buf_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I212 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
pch_25  M31 ( .D(net0203), .B(net0165), .G(dis_pgate_25), .S(net0165));
pch_25  M0 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
pch_25  M9 ( .D(net0166), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
pch_25  M14 ( .D(pump_opamp_out), .B(net125), .G(vref_25), .S(net125));
pch_25  M18 ( .D(net122), .B(vpp_int), .G(net122), .S(vpp_int));
pch_25  M13 ( .D(net124), .B(net125), .G(vdiv), .S(net125));
pch_25  M32 ( .D(dis_pgate_25), .B(vddp_), .G(dis_pgate_25),
     .S(vddp_));
pch_25  M33 ( .D(dis_pgate_25), .B(vddp_), .G(vppdisc_25), .S(vddp_));
pch_25  M12 ( .D(net125), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M19 ( .D(net134), .B(net122), .G(net134), .S(net122));
pch_25  M21 ( .D(net138), .B(net134), .G(net138), .S(net134));
pch_25  M23 ( .D(net142), .B(net138), .G(net142), .S(net138));
pch_25  M24 ( .D(vdiv), .B(net142), .G(vdiv), .S(net142));
pch_25  M25 ( .D(net0224), .B(vdiv), .G(net0224), .S(vdiv));
pch_25  M4_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
pch_25  M4_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
nch_25  M40 ( .D(dis_pgate_25), .B(GND_), .G(vppdisc_25), .S(gnd_));
nch_25  M8 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
nch_25  M16 ( .D(net124), .B(GND_), .G(net124), .S(net155));
nch_25  M17 ( .D(net155), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M6 ( .D(vpp_int), .B(GND_), .G(en_buf_25), .S(net168));
nch_25  M20 ( .D(slow_25), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M7 ( .D(net168), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M41 ( .D(net0224), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M15 ( .D(pump_opamp_out), .B(GND_), .G(net124), .S(net155));
nch_25  M3 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net0250));
rppolywo_m  R5 ( .MINUS(net0165), .PLUS(vpp_int), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(pump_gate), .PLUS(pump_in), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net0247), .PLUS(net0250), .BULK(GND_));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net0247), .BULK(GND_));

endmodule
// Library - NVCM, Cell - ml_vpp_vco, View - schematic
// LAST TIME SAVED: Apr  8 16:31:55 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpp_vco ( clk_25_0, pbias_25, slow_25, en_25, freq_25 );
output  clk_25_0;

inout  pbias_25, slow_25;

input  en_25;

input [1:0]  freq_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:1]  freq_b_25;



nch_na25  M4 ( .D(GND_), .B(GND_), .G(net173), .S(GND_));
nch_na25  M15 ( .D(GND_), .B(GND_), .G(net185), .S(GND_));
nch_na25  M16 ( .D(GND_), .B(GND_), .G(net193), .S(GND_));
nch_na25  M2 ( .D(GND_), .B(GND_), .G(net189), .S(GND_));
nch_25  M5 ( .D(net173), .B(GND_), .G(net185), .S(net177));
nch_25  M6 ( .D(net177), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M13 ( .D(net181), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M14 ( .D(net185), .B(GND_), .G(net193), .S(net181));
nch_25  M8 ( .D(net189), .B(GND_), .G(net173), .S(net201));
nch_25  M17 ( .D(net193), .B(GND_), .G(net195), .S(net197));
nch_25  M18 ( .D(net197), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M1 ( .D(net201), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M23 ( .D(pbias_osc_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M24 ( .D(slow_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M25 ( .D(nbias_osc_25), .B(GND_), .G(en_25), .S(slow_25));
pch_25  M7 ( .D(net173), .B(vddp_), .G(net185), .S(net236));
pch_25  M10 ( .D(net236), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M9 ( .D(net248), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M3 ( .D(net189), .B(vddp_), .G(net173), .S(net248));
pch_25  M11 ( .D(net256), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M12 ( .D(net185), .B(vddp_), .G(net193), .S(net256));
pch_25  M19 ( .D(net193), .B(vddp_), .G(net195), .S(net260));
pch_25  M20 ( .D(net260), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M22 ( .D(pbias_osc_25), .B(vddp_), .G(en_b_25), .S(net228));
pch_25  M26_1_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M26_0_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_1_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_0_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M28 ( .D(net212), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M29 ( .D(nbias_osc_25), .B(vddp_), .G(freq_25[0]), .S(net212));
pch_25  M30 ( .D(nbias_osc_25), .B(vddp_), .G(freq_b_25[1]),
     .S(net208));
pch_25  M21 ( .D(net228), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
nand2_25 I96 ( .G(GND_), .Pb(vddp_), .A(net189), .Y(net195), .P(vddp_),
     .B(en_25), .Gb(GND_));
inv_25 I201 ( .IN(net195), .OUT(clk_25_0), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I188 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I199 ( .IN(freq_25[1]), .OUT(freq_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));

endmodule
// Library - NVCM, Cell - ml_vpp_pump, View - schematic
// LAST TIME SAVED: Apr  7 18:25:20 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpp_pump ( pump_in, clkin_25, en_25 );
inout  pump_in;

input  clkin_25, en_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



// nmoscap_25  C0 ( .MINUS(clk_25), .PLUS(s_0));
// nmoscap_25  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
// nmoscap_25  C7 ( .MINUS(clk_25), .PLUS(s_2));
// nmoscap_25  C1 ( .MINUS(clk_b_25), .PLUS(s_3));
pch_25  M0 ( .D(net23), .B(vddp_), .G(net64), .S(vddp_));
inv_25 I194 ( .IN(clkin_25), .OUT(net70), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(en_25), .OUT(net64), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I210 ( .IN(net28), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I219 ( .IN(net40), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I220 ( .IN(net34), .OUT(net46), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I221 ( .IN(net46), .OUT(net40), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I224 ( .IN(clkin_25), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I209 ( .IN(net70), .OUT(net28), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
nch_na25  M10 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
nch_na25  M11 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
nch_na25  M12 ( .D(s_2), .B(GND_), .G(s_2), .S(s_3));
nch_na25  M22 ( .D(net23), .B(GND_), .G(net23), .S(s_0));
nch_na25  M1 ( .D(s_3), .B(GND_), .G(s_3), .S(pump_in));

endmodule
// Library - NVCM, Cell - ml_vpp_pumpx3, View - schematic
// LAST TIME SAVED: Apr  8 17:28:05 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpp_pumpx3 ( pump_in, clkin_0_25, pumpen_25 );
inout  pump_in;

input  clkin_0_25, pumpen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I195 ( .IN(clkin_0_25), .OUT(net13), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I84 ( .IN(net13), .OUT(net024), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
ml_vpp_pump Ivpp_pump_0 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(clkin_0_25));
ml_vpp_pump I79 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net024));
ml_vpp_pump Ivpp_pump_1 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net13));

endmodule
// Library - NVCM, Cell - ml_vppint_top, View - schematic
// LAST TIME SAVED: Feb 12 09:53:31 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vppint_top ( vpint_en, vpp_int, bgr, fsm_lshven_buf,
     fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf, fsm_pgmvfy_buf,
     fsm_tm_xforce, fsm_tm_xvppint, fsm_vpgmwl_buf, fsm_wgnden_buf );
output  vpint_en;

inout  vpp_int;

input  bgr, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_wgnden_buf;

input [2:0]  fsm_vpgmwl_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_25;

wire  [1:0]  freq_25;



ml_hv2vddp_sw Ivpxa_2vddp_sw ( .hv2vddp(vpp_2_vdd),
     .vddp_tieh(vddp_tieh), .out_hv(vpp_int));
inv_25 I38 ( .IN(vddp_tieh), .OUT(freq_25[1]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I86 ( .IN(vddp_tieh), .OUT(freq_25[0]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
ml_vpp_ref Ivpp_ref ( .vref_25(vref_25), .vppwl_25(vppwl_25[2:0]),
     .pumpen_25(pumpen_25), .bgr(bgr));
ml_vpp_ctrl Ivpp_ctrl ( .vpint_en(vpint_en),
     .fsm_pgmvfy_buf(fsm_pgmvfy_buf), .fsm_nvcmen_buf(fsm_nvcmen_buf),
     .vppdisc_25(vppdisc_25), .fsm_wgnden(fsm_wgnden_buf),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf), .vppwl_25(vppwl_25[2:0]),
     .vpp_2_vdd(vpp_2_vdd), .pumpen_25(pumpen_25));
ml_vpp_reg Ivpp_reg ( .bgr(bgr), .slow_25(slow_25),
     .pbias_25(pbias_25), .vref_25(vref_25), .vppdisc_25(vppdisc_25),
     .pumpen_25(pumpen_25), .pump_in(pump_in), .vpp_int(vpp_int));
ml_vpp_vco Ivpp_vco ( .pbias_25(pbias_25), .slow_25(slow_25),
     .freq_25(freq_25[1:0]), .en_25(pumpen_25), .clk_25_0(clkin_0_25));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));
// nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpp_int));
ml_vpp_pumpx3 Ivpp_pumpx3 ( .pump_in(pump_in), .pumpen_25(pumpen_25),
     .clkin_0_25(clkin_0_25));

endmodule
// Library - NVCM, Cell - UBGR_2511_065_FLAT, View - schematic
// LAST TIME SAVED: Apr  1 15:53:36 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module UBGR_2511_065_FLAT ( VREF, PDN, T0, T1, T2, T3, TEN, VDD25, VSS
     );
output  VREF;

input  PDN, T0, T1, T2, T3, TEN, VDD25, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_bgr_top, View - schematic
// LAST TIME SAVED: Apr  7 14:19:14 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_bgr_top ( bgr_int, fsm_nvcmen_buf, fsm_trim_vbg_buf );
inout  bgr_int;

input  fsm_nvcmen_buf;

input [3:0]  fsm_trim_vbg_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  bgr_trim_25;

wire  [0:3]  net48;

wire  [0:3]  net53;

wire  [0:3]  net44;



inv_25 I38 ( .IN(net58), .OUT(PDN), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
vddp_tiehigh I85 ( .vddp_tieh(TEN));
UBGR_2511_065_FLAT Ibgr ( .TEN(TEN), .VSS(gnd_), .VDD25(vddp_),
     .VREF(bgr_int), .T3(bgr_trim_25[3]), .T2(bgr_trim_25[2]),
     .T1(bgr_trim_25[1]), .T0(bgr_trim_25[0]), .PDN(PDN));
inv_hvt I88_3_ ( .A(fsm_trim_vbg_buf[3]), .Y(net48[0]));
inv_hvt I88_2_ ( .A(fsm_trim_vbg_buf[2]), .Y(net48[1]));
inv_hvt I88_1_ ( .A(fsm_trim_vbg_buf[1]), .Y(net48[2]));
inv_hvt I88_0_ ( .A(fsm_trim_vbg_buf[0]), .Y(net48[3]));
inv_hvt I319 ( .A(net50), .Y(net46));
inv_hvt I87_3_ ( .A(net48[0]), .Y(net44[0]));
inv_hvt I87_2_ ( .A(net48[1]), .Y(net44[1]));
inv_hvt I87_1_ ( .A(net48[2]), .Y(net44[2]));
inv_hvt I87_0_ ( .A(net48[3]), .Y(net44[3]));
inv_hvt I323 ( .A(fsm_nvcmen_buf), .Y(net50));
ml_ls_vdd2vdd25 I80_3_ ( .in(net44[0]), .sup(vddp_),
     .out_vddio_b(net53[0]), .out_vddio(bgr_trim_25[3]),
     .in_b(net48[0]));
ml_ls_vdd2vdd25 I80_2_ ( .in(net44[1]), .sup(vddp_),
     .out_vddio_b(net53[1]), .out_vddio(bgr_trim_25[2]),
     .in_b(net48[1]));
ml_ls_vdd2vdd25 I80_1_ ( .in(net44[2]), .sup(vddp_),
     .out_vddio_b(net53[2]), .out_vddio(bgr_trim_25[1]),
     .in_b(net48[2]));
ml_ls_vdd2vdd25 I80_0_ ( .in(net44[3]), .sup(vddp_),
     .out_vddio_b(net53[3]), .out_vddio(bgr_trim_25[0]),
     .in_b(net48[3]));
ml_ls_vdd2vdd25 I335 ( .in(net46), .sup(vddp_), .out_vddio_b(net58),
     .out_vddio(bgr_en_25), .in_b(net50));

endmodule
// Library - NVCM, Cell - ml_pump_vpxa_3.3v, View - schematic
// LAST TIME SAVED: Feb  6 11:01:23 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_pump_vpxa_3_3v ( out, clkin_25, en );
inout  out;

input  clkin_25, en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M10 ( .B(GND_), .D(s_0), .G(s_0), .S(s_1));
nch_na25  M11 ( .B(GND_), .D(s_1), .G(s_1), .S(s_2));
nch_na25  M12 ( .B(GND_), .D(s_2), .G(s_2), .S(out));
nch_na25  M22 ( .B(GND_), .D(net0115), .G(net0115), .S(s_0));
inv_25 I194 ( .IN(clkin_25), .OUT(net064), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(en), .OUT(net042), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I210 ( .IN(net076), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I219 ( .IN(net040), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I220 ( .IN(net034), .OUT(net046), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I221 ( .IN(net046), .OUT(net040), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I224 ( .IN(clkin_25), .OUT(net034), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I209 ( .IN(net064), .OUT(net076), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
pch_25  M0 ( .D(net0115), .B(vddp_), .G(net042), .S(vddp_));
// nmoscap_25  C0 ( .MINUS(clk_25), .PLUS(s_0));
// nmoscap_25  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
// nmoscap_25  C7 ( .MINUS(clk_25), .PLUS(s_2));

endmodule
// Library - sbtlibn65lp, Cell - ml_dlatch_25, View - schematic
// LAST TIME SAVED: Feb 21 13:49:32 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_dlatch_25 ( Q_25, D_25, EN_25, R_25 );
output  Q_25;

input  D_25, EN_25, R_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M9 ( .D(net31), .B(vddp_), .G(EN_25), .S(vddp_));
pch_25  M7 ( .D(net39), .B(vddp_), .G(EN_B_25), .S(vddp_));
pch_25  M3 ( .D(net52), .B(vddp_), .G(D_25), .S(net39));
pch_25  M4 ( .D(net52), .B(vddp_), .G(Q_25), .S(net31));
nch_25  M8 ( .D(net52), .B(GND_), .G(D_25), .S(net48));
nch_25  M1 ( .D(net48), .B(GND_), .G(EN_25), .S(GND_));
nch_25  M5 ( .D(net40), .B(GND_), .G(EN_B_25), .S(GND_));
nch_25  M6 ( .D(net52), .B(GND_), .G(Q_25), .S(net40));
inv_25 I156 ( .IN(EN_25), .OUT(EN_B_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nor2_25 I161 ( .A(net52), .Y(Q_25), .Gb(GND_), .G(GND_), .Pb(vddp_),
     .P(vddp_), .B(R_25));

endmodule
// Library - NVCM, Cell - ml_pump_clk_reg, View - schematic
// LAST TIME SAVED: Feb 13 16:09:37 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_pump_clk_reg ( clk_out_25, clk_in_25, pump_chrg_25,
     pump_on_25 );
output  clk_out_25;

input  clk_in_25, pump_chrg_25, pump_on_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



exor2_25 I85 ( .A(clk_in_25), .Y(net020), .B(clk_out_25));
nand2_25 I78 ( .G(GND_), .Pb(vddp_), .A(pump_chrg_25), .Y(clk_freeze),
     .P(vddp_), .B(pump_on_25), .Gb(GND_));
inv_25 I72 ( .IN(net020), .OUT(clk_equal), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(vddp_tieh), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
vddp_tiehigh I117 ( .vddp_tieh(vddp_tieh));
ml_dlatch_25 I63 ( .D_25(clk_in_25), .EN_25(clk_go), .R_25(net34),
     .Q_25(clk_out_25));
ml_dlatch_25 I64 ( .D_25(vddp_tieh), .EN_25(clk_equal),
     .R_25(clk_freeze), .Q_25(clk_go));

endmodule
// Library - misc, Cell - vpp_clamp, View - schematic
// LAST TIME SAVED: May  1 10:47:24 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module vpp_clamp ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



vpp_clamp_finger I0_9_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_8_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_7_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_6_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_5_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_4_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_3_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_2_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_1_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_0_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));

endmodule
// Library - NVCM, Cell - ml_pump_vpxa_x2, View - schematic
// LAST TIME SAVED: Feb  6 11:01:27 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_pump_vpxa_x2 ( vpxa_int, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, pumpen, pumpen_25, vpxa_clk_25, vpxa_clk_b_25 );
inout  vpxa_int;

input  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25, pumpen,
     pumpen_25, vpxa_clk_25, vpxa_clk_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_pump_vpxa_3_3v Ivpxa_pump_0 ( .en(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_0_25));
ml_pump_vpxa_3_3v Ivpxa_pump_2 ( .en(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_2_25));
ml_pump_vpxa_3_3v Ivpxa_pump_1 ( .en(pumpen_25), .clkin_25(clkin_1_25),
     .out(vpxa_int));
ml_pump_clk_reg Iclk_reg_0 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_0_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_0_25));
ml_pump_clk_reg Iclk_reg_2 ( .clk_in_25(vpxa_clk_b_25),
     .pump_chrg_25(pump_chrg_2_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_2_25));
ml_pump_clk_reg Iclk_reg_1 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_1_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_1_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_osc, View - schematic
// LAST TIME SAVED: Mar 14 15:11:03 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpxa_osc ( vpxa_clk_25, bgr, freq_25, pumpen_25 );
output  vpxa_clk_25;

inout  bgr;

input  pumpen_25;

input [1:0]  freq_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  freq_buf_b_25;



inv_25 I38 ( .IN(pumpen_25), .OUT(pbiasen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I195 ( .IN(freq_25[0]), .OUT(freq_buf_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
pch_25  M9 ( .D(net64), .B(vddp_), .G(pbiasen_b_25), .S(vddp_));
pch_25  M4_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
pch_25  M4_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
pch_25  M0 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
nch_25  M8 ( .D(pbias_25), .B(GND_), .G(pbiasen_b_25), .S(gnd_));
nch_25  M3 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net74));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net83), .PLUS(net74), .BULK(GND_));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net83), .BULK(GND_));
ml_vpp_vco Ivpx_vpp_vco ( .pbias_25(pbias_25), .slow_25(net86),
     .freq_25({freq_25[1], freq_buf_b_25[0]}), .en_25(pumpen_25),
     .clk_25_0(vpxa_clk_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_ctrl, View - schematic
// LAST TIME SAVED: Feb  6 11:01:40 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpxa_ctrl ( pumpen, pumpen_25, vpxa_2_vdd, fsm_pumpen,
     fsm_tm_xforce, fsm_tm_xvpxaint );
output  pumpen, pumpen_25, vpxa_2_vdd;

input  fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I73 ( .A(fsm_tm_xvpxaint), .B(fsm_tm_xforce), .Y(net042));
inv_25 I38 ( .IN(net045), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I173 ( .in(net049), .sup(vddp_), .out_vddio_b(net045),
     .out_vddio(net046), .in_b(net075));
nor2_hvt I72 ( .A(vpxa_off), .B(net065), .Y(net049));
nor2_hvt I69 ( .A(vpxa_2_vdd), .B(vpxa_2_vdd), .Y(net043));
inv_hvt I75 ( .A(net049), .Y(net056));
inv_hvt I76 ( .A(net056), .Y(pumpen));
inv_hvt I110 ( .A(net049), .Y(net075));
inv_hvt I74 ( .A(net042), .Y(net065));
inv_hvt I131 ( .A(fsm_pumpen), .Y(vpxa_2_vdd));
inv_hvt I70 ( .A(net043), .Y(vpxa_off));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff_25, View - schematic
// LAST TIME SAVED: Feb 11 11:37:05 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_dff_25 ( Q_25, Q_B_25, CLK_25, D_25, R_25 );
output  Q_25, Q_B_25;

input  CLK_25, D_25, R_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I87 ( .IN(net044), .OUT(net038), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I72 ( .IN(CLK_25), .OUT(net044), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I90 ( .IN(Q_25), .OUT(Q_B_25), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
ml_dlatch_25 Ilatch2 ( .D_25(net053), .EN_25(net038), .R_25(R_25),
     .Q_25(Q_25));
ml_dlatch_25 Ilatch1 ( .Q_25(net053), .EN_25(net044), .D_25(D_25),
     .R_25(R_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp_n, View - schematic
// LAST TIME SAVED: Feb  5 15:08:44 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_core_sa_comp_n ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M0 ( .D(out_div), .B(vddp_), .G(out_ref), .S(vddp_));
pch_25  M4 ( .D(out_ref), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M5 ( .D(out_div), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M7 ( .D(out_ref), .B(vddp_), .G(out_ref), .S(vddp_));
nch_25  M1 ( .D(out_div), .B(GND_), .G(in_div), .S(net049));
nch_25  M2 ( .D(out_ref), .B(GND_), .G(in_ref), .S(net049));
nch_25  M6_1_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp_top_n, View - schematic
// LAST TIME SAVED: Feb 21 13:55:00 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_core_sa_comp_top_n ( pump_chrg_25, in_div, in_ref, sa_bias,
     saen_25 );
output  pump_chrg_25;

input  in_div, in_ref, sa_bias, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_25 I103 ( .G(gnd_), .Pb(vddp_), .A(saen_25), .Y(chrg_b_25),
     .P(vddp_), .B(net27), .Gb(gnd_));
nch_25  M6_1_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
inv_25 I102 ( .IN(chrg_b_25), .OUT(pump_chrg_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I104 ( .IN(out_div2), .OUT(net27), .P(vddp_), .Pb(vddp_),
     .G(net087), .Gb(gnd_));
ml_core_sa_comp_n Icore_sa_comp_n0 ( .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp_n Iml_core_sa_comp_n1 ( .out_div(out_div2),
     .out_ref(out_ref2), .in_div(in_div2), .in_ref(in_ref2),
     .sa_bias(sa_bias), .saen_25(saen_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_reg, View - schematic
// LAST TIME SAVED: May  3 13:50:36 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpxa_reg ( freq_25, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, vpxa_int, bgr, fsm_vrdwl, pumpen, vpxa_clk_25 );
output  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25;

inout  vpxa_int;

input  bgr, pumpen, vpxa_clk_25;

output [1:0]  freq_25;

input [2:0]  fsm_vrdwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  freq_in_25;

wire  [0:2]  vrdwl_vpxa;

wire  [0:2]  vrdwl_b_vpxa;



nand2_25 I145 ( .G(GND_), .Pb(vddp_), .A(net0171), .Y(freq_in_25[0]),
     .P(vddp_), .B(net0179), .Gb(GND_));
nand2_25 I158 ( .G(GND_), .Pb(vddp_), .A(net0179), .Y(freq_in_25[1]),
     .P(vddp_), .B(net0163), .Gb(GND_));
nand3_25 I44 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0179),
     .C(pump_chrg_0_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I149 ( .B(pump_chrg_1_b_25), .A(pump_chrg_2_25), .Y(net0171),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I159 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0163),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
ml_dff_25 I125 ( .Q_B_25(net0187), .R_25(saen_b_25),
     .D_25(freq_in_25[1]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[1]));
ml_dff_25 I126 ( .Q_B_25(net0192), .R_25(saen_b_25),
     .D_25(freq_in_25[0]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[0]));
inv_hvt I85 ( .A(net171), .Y(net175));
inv_hvt I183 ( .A(fsm_vrdwl[2]), .Y(net171));
inv_hvt I83 ( .A(pumpen), .Y(net143));
inv_hvt I82 ( .A(net143), .Y(net145));
inv_hvt I184 ( .A(fsm_vrdwl[1]), .Y(net176));
inv_hvt I187 ( .A(fsm_vrdwl[0]), .Y(net181));
inv_hvt I186 ( .A(net181), .Y(net185));
inv_hvt I185 ( .A(net176), .Y(net180));
inv_25 I155 ( .IN(pump_chrg_0_25), .OUT(pump_chrg_0_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
inv_25 I63 ( .IN(net169), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(net168), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I154 ( .IN(pump_chrg_1_25), .OUT(pump_chrg_1_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_ls_vdd2vdd25 I191 ( .in(saen_25), .sup(vpxa_int),
     .out_vddio_b(saen_b_vpxa), .out_vddio(net0210), .in_b(saen_b_25));
ml_ls_vdd2vdd25 I335 ( .in(net145), .sup(vddp_), .out_vddio_b(net168),
     .out_vddio(net169), .in_b(net143));
ml_ls_vdd2vdd25 I87 ( .in(net171), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[2]), .out_vddio(vrdwl_b_vpxa[2]),
     .in_b(net175));
ml_ls_vdd2vdd25 I98 ( .in(net176), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[1]), .out_vddio(vrdwl_b_vpxa[1]),
     .in_b(net180));
ml_ls_vdd2vdd25 I99 ( .in(net181), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[0]), .out_vddio(vrdwl_b_vpxa[0]),
     .in_b(net185));
ml_core_sa_comp_top_n Icore_sa_comp_top_n2 (
     .pump_chrg_25(pump_chrg_2_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_2));
ml_core_sa_comp_top_n core_sa_comp_top_n0 (
     .pump_chrg_25(pump_chrg_0_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_0));
ml_core_sa_comp_top_n Icore_sa_comp_top_n1 (
     .pump_chrg_25(pump_chrg_1_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_1));
rppolywo_m  R29 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R28 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R20 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R27 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(in_div_0), .PLUS(net202), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net232), .PLUS(net223), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(net270), .PLUS(net226), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net226), .PLUS(net229), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(sa_bias), .PLUS(net232), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net202), .PLUS(net237), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(net237), .PLUS(net270), .BULK(GND_));
rppolywo_m  R30 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(gnd_), .PLUS(in_div_2), .BULK(GND_));
rppolywo_m  R31 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
pch_25  M3 ( .D(net229), .B(vpxa_int), .G(saen_b_vpxa), .S(vpxa_int));
pch_25  M11_1_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M11_0_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M15 ( .D(net237), .B(vpxa_int), .G(vrdwl_vpxa[0]), .S(net270));
pch_25  M37 ( .D(net226), .B(vpxa_int), .G(vrdwl_vpxa[2]), .S(net229));
pch_25  M1 ( .D(net223), .B(vddp_), .G(saen_b_25), .S(vddp_));
pch_25  M14 ( .D(net270), .B(vpxa_int), .G(vrdwl_vpxa[1]), .S(net226));
pch_25  M8_1_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
pch_25  M8_0_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
nch_25  M2 ( .D(sa_bias), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M32 ( .D(net229), .B(GND_), .G(vrdwl_b_vpxa[2]), .S(net226));
nch_25  M0_3_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_2_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_1_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_0_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M9 ( .D(net270), .B(GND_), .G(vrdwl_b_vpxa[0]), .S(net237));
nch_25  M7 ( .D(net226), .B(GND_), .G(vrdwl_b_vpxa[1]), .S(net270));

endmodule
// Library - NVCM, Cell - ml_hv2vdd_sw, View - schematic
// LAST TIME SAVED: Apr  8 14:27:39 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_hv2vdd_sw ( out_hv, hv2vdd, vddp_tieh );
inout  out_hv;

input  hv2vdd, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M1 ( .D(net27), .B(GND_), .G(vddp_tieh), .S(out_hv));
nch_na25  M2 ( .D(vdd_), .B(GND_), .G(hv2vdd_25), .S(net27));
inv_25 I62 ( .IN(net40), .OUT(hv2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net40),
     .out_vddio(net37), .in_b(net46));
inv_hvt I65 ( .A(hv2vdd), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));

endmodule
// Library - NVCM, Cell - ml_vpxa_top, View - schematic
// LAST TIME SAVED: Sep  3 10:36:27 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_vpxa_top ( vpxa_int, bgr, fsm_pumpen, fsm_tm_xforce,
     fsm_tm_xvpxaint, fsm_vrdwl );
inout  vpxa_int;

input  bgr, fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;

input [2:0]  fsm_vrdwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  freq_25;



// nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpxa_int));
ml_pump_vpxa_x2 Ipump_vpxa_x3 ( .pumpen(pumpen),
     .vpxa_clk_b_25(vpxa_clk_b_25), .vpxa_clk_25(vpxa_clk_25),
     .pumpen_25(pumpen_25), .pump_chrg_2_25(pump_chrg_2_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_0_25(pump_chrg_0_25),
     .vpxa_int(vpxa_int));
inv_25 I73 ( .IN(vpxa_clk_25), .OUT(vpxa_clk_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_vpxa_osc Ivpxa_osc ( .freq_25(freq_25[1:0]), .bgr(bgr),
     .pumpen_25(pumpen_25), .vpxa_clk_25(vpxa_clk_25));
ml_vpxa_ctrl Ivpxa_ctrl ( .fsm_pumpen(fsm_pumpen), .pumpen(pumpen),
     .pumpen_25(pumpen_25), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .vpxa_2_vdd(vpxa_2_vdd));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));
ml_vpxa_reg Ivpxa_reg ( .pump_chrg_0_25(pump_chrg_0_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_2_25(pump_chrg_2_25),
     .freq_25(freq_25[1:0]), .vpxa_clk_25(vpxa_clk_25),
     .pumpen(pumpen), .fsm_vrdwl(fsm_vrdwl[2:0]), .bgr(bgr),
     .vpxa_int(vpxa_int));
ml_hv2vdd_sw Ivpxa_2vdd_sw ( .vddp_tieh(vddp_tieh),
     .hv2vdd(vpxa_2_vdd), .out_hv(vpxa_int));

endmodule
// Library - NVCM, Cell - ml_hvmux_top_ctrl, View - schematic
// LAST TIME SAVED: May  2 18:30:47 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_hvmux_top_ctrl ( bgrext_en, bgrint_en, en_vblinhi,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp, fsm_lshven,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint, fsm_wgnden,
     fsm_wpen, tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );
output  bgrext_en, bgrint_en, en_vblinhi, ngate_vddp, ngate_vpxa,
     sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint,
     vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint, vpxaint_ext,
     vtmode, ysup25_2vdd, ysup25_2vddp;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_testdec,
     tm_wleqbl, vpint_en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



mux2_hvt I260 ( .in1(fsm_wgnden), .in0(fsm_wpen), .out(net0217),
     .sel(pgmpulse_b));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
anor21_hvt I245 ( .A(net0189), .B(net0193), .Y(vppint_ext),
     .C(net0188));
anor21_hvt I109 ( .A(net0201), .B(net0199), .Y(vpxa_ext), .C(net0188));
nand3_hvt I248 ( .Y(net0189), .B(vpint_en), .C(fsm_tm_xvppint),
     .A(fsm_tm_xforce));
nand3_hvt I246 ( .Y(net0201), .B(vddp_rd_b), .C(fsm_tm_xvpxa),
     .A(fsm_tm_xforce));
nand3_hvt I247 ( .Y(net0193), .B(pmprd), .C(pmprd),
     .A(fsm_tm_xvppint));
nand3_hvt I35 ( .C(fsm_lshven), .A(fsm_pgm), .Y(pgmpulse_b),
     .B(net0327));
nand3_hvt I205 ( .Y(net0213), .B(net0321), .C(pgmpulse_b),
     .A(net0321));
nand3_hvt I240 ( .C(pmprd), .A(fsm_tm_xvpxa), .Y(net0199), .B(pmprd));
nor2_hvt I213 ( .A(net0324), .B(fsm_nvcmen_b), .Y(net0251));
nor2_hvt I224 ( .A(vddp_rd_b), .B(net0258), .Y(vpxa_vppd));
nor2_hvt I214 ( .A(net0251), .B(net0266), .Y(sbhvsup_vppint));
nor2_hvt I215 ( .A(net0264), .B(net0311), .Y(sbhvsup_vddp));
nor2_hvt I183 ( .A(net87), .B(net73), .Y(ysup25_2vddp));
nor2_hvt I14 ( .A(net75), .B(net93), .Y(ysup25_2vdd));
nor2_hvt I207 ( .A(net0325), .B(net0260), .Y(sb25sup_vddp));
nor2_hvt I206 ( .A(net0268), .B(net0213), .Y(sb25sup_vpxa));
nor2_hvt I185 ( .A(gnd_tiel), .B(gnd_tiel), .Y(net0240));
nor2_hvt I223 ( .B(net0240), .Y(vddp_rd), .A(net0349));
nor2_hvt I195 ( .A(net0272), .B(rd_vddp), .Y(ngate_vpxa));
nor2_hvt I196 ( .A(net0331), .B(net0270), .Y(ngate_vddp));
nor2_hvt I225 ( .A(net0256), .B(vddp_rd), .Y(vpxa_vpxaint));
ml_pump_a_clkdly I219 ( .in(ysup25_2vddp_b), .out(net75));
ml_pump_a_clkdly I227 ( .in(net0297), .out(net0256));
ml_pump_a_clkdly I226 ( .in(net0319), .out(net0258));
ml_pump_a_clkdly I209 ( .in(net0323), .out(net0260));
ml_pump_a_clkdly I184 ( .in(ysup25_2vdd_b), .out(net73));
ml_pump_a_clkdly I217 ( .in(net0313), .out(net0264));
ml_pump_a_clkdly I216 ( .in(net0309), .out(net0266));
ml_pump_a_clkdly I208 ( .in(net0329), .out(net0268));
ml_pump_a_clkdly I198 ( .in(net0339), .out(net0270));
ml_pump_a_clkdly I197 ( .in(net0335), .out(net0272));
nand2_hvt I254 ( .A(bgrext_en), .Y(bgrint_en), .B(fsm_tm_xforce));
nand2_hvt I104 ( .A(fsm_nvcmen), .Y(net77), .B(tm_wleqbl));
nand2_hvt I179 ( .A(fsm_nvcmen), .Y(net80), .B(net0217));
nand2_hvt I252 ( .A(fsm_nvcmen_buf), .Y(net0277), .B(fsm_tm_xvbg));
nand2_hvt I234 ( .A(fsm_pumpen), .Y(net0286), .B(fsm_tm_xvpxaint));
inv_hvt I259 ( .A(pgmpulse_b), .Y(net0324));
inv_hvt I229 ( .A(vpxa_vppd), .Y(net0297));
inv_hvt I250 ( .A(fsm_pumpen), .Y(net0188));
inv_hvt I182 ( .A(ysup25_2vdd), .Y(ysup25_2vdd_b));
inv_hvt I230 ( .A(vddp_rd), .Y(vddp_rd_b));
inv_hvt I249 ( .A(pgmpulse_b), .Y(pgmpulse));
inv_hvt I131 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I178 ( .A(net77), .Y(vtmode));
inv_hvt I180 ( .A(net80), .Y(net93));
inv_hvt I253 ( .A(net0277), .Y(bgrext_en));
inv_hvt I218 ( .A(sbhvsup_vddp), .Y(net0309));
inv_hvt I221 ( .A(net0251), .Y(net0311));
inv_hvt I220 ( .A(sbhvsup_vppint), .Y(net0313));
inv_hvt I134 ( .A(net93), .Y(net87));
inv_hvt I181 ( .A(ysup25_2vddp), .Y(ysup25_2vddp_b));
inv_hvt I228 ( .A(vpxa_vpxaint), .Y(net0319));
inv_hvt I204 ( .A(rd_vddp), .Y(net0321));
inv_hvt I212 ( .A(sb25sup_vpxa), .Y(net0323));
inv_hvt I210 ( .A(net0213), .Y(net0325));
inv_hvt I202 ( .A(fsm_pgmvfy), .Y(net0327));
inv_hvt I211 ( .A(sb25sup_vddp), .Y(net0329));
inv_hvt I199 ( .A(rd_vddp), .Y(net0331));
inv_hvt I236 ( .A(fsm_tm_xforce), .Y(pmprd));
inv_hvt I200 ( .A(ngate_vddp), .Y(net0335));
inv_hvt I235 ( .A(net0286), .Y(vpxaint_ext));
inv_hvt I201 ( .A(ngate_vpxa), .Y(net0339));
inv_hvt I233 ( .A(fsm_nvcmen_b), .Y(fsm_nvcmen_buf));
nor3_hvt I105 ( .B(tm_testdec), .Y(en_vblinhi), .A(fsm_nvcmen_b),
     .C(tm_allbl_l));
nor3_hvt I186 ( .C(fsm_rd), .A(fsm_tm_rd_mode), .B(fsm_pgmvfy),
     .Y(net0349));
nor3_hvt I187 ( .B(net0240), .Y(rd_vddp), .A(net0349),
     .C(fsm_nvcmen_b));

endmodule
// Library - io, Cell - pvpp, View - schematic
// LAST TIME SAVED: May  1 10:46:55 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module pvpp ( vpp, vppin );
inout  vpp, vppin;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo_m  R1 ( .MINUS(vpp), .PLUS(vppin), .BULK(gnd_));
vddp_tiehigh I60_7_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_6_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_5_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_4_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_3_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_2_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_1_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_0_ ( .vddp_tieh(vddio_in));
vpp_clamp I59_3_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_2_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_1_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_0_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));

endmodule
// Library - NVCM, Cell - ml_hvmux_ls25, View - schematic
// LAST TIME SAVED: Feb 15 14:23:11 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_hvmux_ls25 ( bgrext_en_25, bgrint_en_25, ngate_vddp_25,
     ngate_vpxa_25, sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25, bgrext_en, bgrint_en,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp );
output  bgrext_en_25, bgrint_en_25, ngate_vddp_25, ngate_vpxa_25,
     sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25;

input  bgrext_en, bgrint_en, ngate_vddp, ngate_vpxa, sb25sup_vddp,
     sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint, vppint_ext, vpxa_ext,
     vpxa_vppd, vpxa_vpxaint, vpxaint_ext, vtmode, ysup25_2vdd,
     ysup25_2vddp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I317 ( .A(net054), .Y(net052));
inv_hvt I314 ( .A(vpxa_vppd), .Y(net054));
inv_hvt I327 ( .A(net066), .Y(net056));
inv_hvt I329 ( .A(bgrint_en), .Y(net058));
inv_hvt I321 ( .A(vpxaint_ext), .Y(net060));
inv_hvt I320 ( .A(net060), .Y(net062));
inv_hvt I325 ( .A(net082), .Y(net064));
inv_hvt I326 ( .A(vppint_ext), .Y(net066));
inv_hvt I312 ( .A(bgrext_en), .Y(net068));
inv_hvt I313 ( .A(net068), .Y(net070));
inv_hvt I328 ( .A(net058), .Y(net0487));
inv_hvt I239 ( .A(sb25sup_vpxa), .Y(net0486));
inv_hvt I319 ( .A(net0112), .Y(net0488));
inv_hvt I240 ( .A(net0486), .Y(net080));
inv_hvt I324 ( .A(vpxa_ext), .Y(net082));
inv_hvt I206 ( .A(vtmode), .Y(net084));
inv_hvt I213 ( .A(ysup25_2vdd), .Y(net086));
inv_hvt I214 ( .A(net086), .Y(net088));
inv_hvt I205 ( .A(net084), .Y(net090));
inv_hvt I216 ( .A(net088), .Y(net092));
inv_hvt I110 ( .A(net072), .Y(net074));
inv_hvt I227 ( .A(net098), .Y(net096));
inv_hvt I228 ( .A(ngate_vddp), .Y(net098));
inv_hvt I217 ( .A(net092), .Y(ysup25_2vdd_buf));
inv_hvt I190 ( .A(ysup25_2vddp), .Y(net072));
inv_hvt I219 ( .A(ngate_vpxa), .Y(net0104));
inv_hvt I220 ( .A(net0104), .Y(net0106));
inv_hvt I232 ( .A(sb25sup_vddp), .Y(net0108));
inv_hvt I231 ( .A(net0108), .Y(net0110));
inv_hvt I323 ( .A(vpxa_vpxaint), .Y(net0112));
inv_hvt I256 ( .A(net0116), .Y(net0114));
inv_hvt I257 ( .A(sbhvsup_vddp), .Y(net0116));
inv_hvt I258 ( .A(net0120), .Y(net0118));
inv_hvt I259 ( .A(sbhvsup_vppint), .Y(net0120));
ml_ls_vdd2vdd25 I336 ( .in(net064), .sup(vddp_), .out_vddio_b(net0123),
     .out_vddio(net0207), .in_b(net082));
ml_ls_vdd2vdd25 I337 ( .in(net056), .sup(vddp_), .out_vddio_b(net0128),
     .out_vddio(net0208), .in_b(net066));
ml_ls_vdd2vdd25 I338 ( .in(net052), .sup(vddp_), .out_vddio_b(net0133),
     .out_vddio(net0211), .in_b(net054));
ml_ls_vdd2vdd25 I339 ( .in(net0487), .sup(vddp_),
     .out_vddio_b(net0138), .out_vddio(net0209), .in_b(net058));
ml_ls_vdd2vdd25 I332 ( .in(net070), .sup(vddp_), .out_vddio_b(net0148),
     .out_vddio(net0149), .in_b(net068));
ml_ls_vdd2vdd25 I238 ( .in(net080), .sup(vddp_), .out_vddio_b(net0153),
     .out_vddio(net0154), .in_b(net0486));
ml_ls_vdd2vdd25 I334 ( .in(net062), .sup(vddp_), .out_vddio_b(net0158),
     .out_vddio(net0214), .in_b(net060));
ml_ls_vdd2vdd25 I335 ( .in(net0488), .sup(vddp_),
     .out_vddio_b(net0163), .out_vddio(net0206), .in_b(net0112));
ml_ls_vdd2vdd25 I212 ( .in(net088), .sup(vddp_), .out_vddio_b(net0168),
     .out_vddio(net0169), .in_b(net086));
ml_ls_vdd2vdd25 I226 ( .in(net096), .sup(vddp_), .out_vddio_b(net0173),
     .out_vddio(net0174), .in_b(net098));
ml_ls_vdd2vdd25 I203 ( .in(net072), .sup(vddp_), .out_vddio_b(net077),
     .out_vddio(net078), .in_b(net074));
ml_ls_vdd2vdd25 I221 ( .in(net0106), .sup(vddp_),
     .out_vddio_b(net0183), .out_vddio(net0184), .in_b(net0104));
ml_ls_vdd2vdd25 I233 ( .in(net0110), .sup(vddp_),
     .out_vddio_b(net0188), .out_vddio(net0219), .in_b(net0108));
ml_ls_vdd2vdd25 I207 ( .in(net090), .sup(vddp_), .out_vddio_b(net0193),
     .out_vddio(net0194), .in_b(net084));
ml_ls_vdd2vdd25 I260 ( .in(net0114), .sup(vddp_),
     .out_vddio_b(net0198), .out_vddio(net0220), .in_b(net0116));
ml_ls_vdd2vdd25 I261 ( .in(net0118), .sup(vddp_),
     .out_vddio_b(net0203), .out_vddio(net0204), .in_b(net0120));
inv_25 I390 ( .IN(net0148), .OUT(bgrext_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I384 ( .IN(net0163), .OUT(vpxa_vpxaint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I386 ( .IN(net0133), .OUT(vpxa_vppd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I388 ( .IN(net0123), .OUT(vpxa_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I376 ( .IN(net0168), .OUT(ysup25_2vdd_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I387 ( .IN(net0158), .OUT(vpxaint_ext_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I389 ( .IN(net0128), .OUT(vppint_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I362 ( .IN(net077), .OUT(ysup25_2vddp_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I383 ( .IN(net0203), .OUT(sbhvsup_vppint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I379 ( .IN(net0183), .OUT(ngate_vpxa_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I377 ( .IN(net0193), .OUT(vtmode_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I378 ( .IN(net0173), .OUT(ngate_vddp_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I381 ( .IN(net0153), .OUT(sb25sup_vpxa_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I382 ( .IN(net0198), .OUT(sbhvsup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I380 ( .IN(net0188), .OUT(sb25sup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I391 ( .IN(net0138), .OUT(bgrint_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_bgrxcvr, View - schematic
// LAST TIME SAVED: Apr  8 10:30:41 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_hvmux_bgrxcvr ( bgr, bgr_int, bgrint_en_25, vpp,
     bgrext_en_25, vddp_tieh );
inout  bgr, bgr_int, bgrint_en_25, vpp;

input  bgrext_en_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M0 ( .D(bgr), .B(GND_), .G(bgrint_en_25), .S(bgr_int));
nch_25  M2 ( .D(vpp), .B(GND_), .G(vddp_tieh), .S(net53));
nch_25  M3 ( .D(net53), .B(GND_), .G(bgrext_en_25), .S(bgr));

endmodule
// Library - NVCM, Cell - ml_ysup_25_switch, View - schematic
// LAST TIME SAVED: Apr  8 10:33:54 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_ysup_25_switch ( vdd, vddp, ysup_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25 );
inout  vdd, vddp, ysup_25;

input  ysup25_2vdd_25, ysup25_2vdd_buf, ysup25_2vddp_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd), .B(GND_), .G(ysup25_2vdd_25), .S(ysup_25));
pch_25  M5 ( .D(net73), .B(vddp), .G(ysup25_2vddp_b_25), .S(vddp));
pch_25  M0 ( .D(ysup_25), .B(ysup_25), .G(ysup25_2vdd_buf), .S(net73));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_vblinhi, View - schematic
// LAST TIME SAVED: Feb  1 08:51:27 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_ymux_ctrl_vblinhi ( vblinhi, vpxa, en_vblinhi, vtmode,
     vtmode_25 );
inout  vblinhi, vpxa;

input  en_vblinhi, vtmode, vtmode_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I191 ( .A(en_vblinhi), .B(vtmode_buf), .Y(ngate_inhi_lv));
nand2_hvt I104 ( .A(net063), .Y(pgate_inhi_lv), .B(en_vblinhi));
inv_hvt I110 ( .A(net063), .Y(vtmode_buf));
inv_hvt I190 ( .A(vtmode), .Y(net063));
nch_25  M9 ( .D(net062), .B(GND_), .G(net062), .S(vblinhi));
nch_25  M8 ( .D(vpxa), .B(GND_), .G(vtmode_25), .S(net062));
pch_hvt  M7_1_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_0_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
nch_hvt  M0_1_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_0_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_top, View - schematic
// LAST TIME SAVED: May  2 18:49:30 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_hvmux_top ( bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi, vpp, vpp_int, vpxa, vpxa_int, ysup_25, fsm_lshven,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint, fsm_wgnden,
     fsm_wpen, tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );
inout  bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi, vpp,
     vpp_int, vpxa, vpxa_int, ysup_25;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_testdec,
     tm_wleqbl, vpint_en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ixcvr_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(vppint_ext_25), .hv_in_hv(vpp_int), .hv_out_hv(vpp));
ml_hvmux_top_ctrl Ihvmux_top_ctrl ( .vpint_en(vpint_en),
     .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl),
     .tm_testdec(tm_testdec), .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvpxa(fsm_tm_xvpxa), .fsm_tm_xvppint(fsm_tm_xvppint),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .ysup25_2vddp(ysup25_2vddp), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vppint(sbhvsup_vppint), .sbhvsup_vddp(sbhvsup_vddp),
     .sb25sup_vpxa(sb25sup_vpxa), .sb25sup_vddp(sb25sup_vddp),
     .ngate_vpxa(ngate_vpxa), .ngate_vddp(ngate_vddp),
     .en_vblinhi(en_vblinhi), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en));
ml_hvmux_ls25 Ihvmux_ls25 ( .ysup25_2vddp(ysup25_2vddp),
     .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vppint_25(sbhvsup_vppint_25), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en), .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vtmode_25(vtmode_25),
     .vpxaint_ext_25(vpxaint_ext_25),
     .vpxa_vpxaint_25(vpxa_vpxaint_25), .vpxa_vppd_25(vpxa_vppd_25),
     .vpxa_ext_25(net164), .vppint_ext_25(vppint_ext_25),
     .sbhvsup_vddp_25(sbhvsup_vddp_25),
     .sb25sup_vpxa_25(sb25sup_vpxa_25),
     .sb25sup_vddp_25(sb25sup_vddp_25), .ngate_vpxa_25(ngate_vpxa_25),
     .ngate_vddp_25(ngate_vddp_25), .bgrint_en_25(bgrint_en_25),
     .bgrext_en_25(bgrext_en_25));
ml_hvmux_bgrxcvr Ixcvr_bgr ( .vddp_tieh(vddp_tieh),
     .bgrext_en_25(bgrext_en_25), .vpp(vpp),
     .bgrint_en_25(bgrint_en_25), .bgr_int(bgr_int), .bgr(bgr));
ml_hv_hotswitch Ixcvr_vpxa_int ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa_int), .hv_out_hv(vpp));
ml_hv_hotswitch Ixcvr_vpxa ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa), .hv_out_hv(vpp));
ml_hvmux_hotswitch Isw_sbhvsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(sbhvsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sb25sup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sb25sup_vpxa_25), .sel_hv_a_25(sb25sup_vddp_25),
     .out_hv(sb25sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_ngate ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(ngate_vpxa_25), .sel_hv_a_25(ngate_vddp_25),
     .out_hv(ngate_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_1_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vpxa_int), .hvin_a_hv(vpxa_int));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_0_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vpxa_int), .hvin_a_hv(vpxa_int));
ml_ysup_25_switch Isw_ysup25_1_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ysup_25_switch Isw_ysup25_0_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
vddp_tiehigh I188_9_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_8_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_0_ ( .vddp_tieh(vddp_tieh));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_1_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_0_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));

endmodule
// Library - NVCM, Cell - ml_chip_nvcm_1f, View - schematic
// LAST TIME SAVED: Feb 17 11:56:19 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_chip_nvcm_1f ( nv_dataout, vpp, fsm_blkadd, fsm_blkadd_b,
     fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_trim_vbg,
     fsm_vpgmwl, fsm_vpxaset, fsm_vrdwl, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbl_h, tm_allbl_l, tm_allwl_h,
     tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr, tm_wleqbl );

inout  vpp;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint,
     fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr, tm_wleqbl;

output [8:0]  nv_dataout;

input [3:0]  fsm_trim_ipp;
input [3:0]  fsm_blkadd;
input [7:0]  fsm_rowadd;
input [3:0]  fsm_trim_vbg;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefpgm;
input [2:0]  fsm_vrdwl;
input [3:0]  fsm_blkadd_b;
input [2:0]  fsm_vpgmwl;
input [2:0]  fsm_trim_rrefrd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  fsm_trim_vbg_buf;

wire  [2:0]  fsm_vpgmwl_buf;



ml_chip_spare Ich_spare_2 ( );
ml_core_1f Icore_1f ( .fsm_pgmdisc(fsm_pgmdisc), .fsm_din(fsm_din),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol), .tm_dma(tm_dma),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_nv_bstream(fsm_nv_bstream),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_blkadd(fsm_blkadd[3:0]), .bgr(bgr), .ngate_25(ngate_25),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpp_int(vpp_int),
     .vpxa(vpxa), .ysup_25(ysup_25), .nv_dataout(nv_dataout[8:0]),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));
// nmoscap_25  C7 ( .MINUS(GND_), .PLUS(vddp_));
// nmoscap_25  C0 ( .MINUS(GND_), .PLUS(vpxa));
ml_chip_buf_top Ichip_buf_top ( .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmvfy_buf(fsm_pgmvfy_buf), .fsm_pgm(fsm_pgm),
     .fsm_pgm_buf(fsm_pgm_buf), .fsm_wgnden_buf(fsm_wgnden_buf),
     .fsm_wgnden(fsm_wgnden), .fsm_vpgmwl(fsm_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_nvcmen(fsm_nvcmen), .fsm_lshven(fsm_lshven),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .fsm_lshven_buf(fsm_lshven_buf));
ml_vppint_top Ivppint_top ( .vpint_en(vpint_en),
     .fsm_pgmvfy_buf(fsm_pgmvfy_buf), .fsm_nvcmen_buf(fsm_nvcmen_buf),
     .vpp_int(vpp_int), .fsm_wgnden_buf(fsm_wgnden_buf), .bgr(bgr),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf));
ml_bgr_top Ibgr_top ( .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .bgr_int(bgr_int));
ml_vpxa_top Ivpxa_top ( .fsm_pumpen(fsm_pumpen),
     .fsm_vrdwl(fsm_vrdwl[2:0]), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .bgr(bgr), .vpxa_int(vpxa));
ml_hvmux_top Ihvmux_top ( .vpint_en(vpint_en), .fsm_wpen(fsm_wpen),
     .tm_wleqbl(tm_wleqbl), .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden_buf), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvpxa(fsm_tm_xvpxa), .fsm_tm_xvppint(fsm_tm_xvppint),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy_buf),
     .fsm_pgm(fsm_pgm_buf), .fsm_nvcmen(fsm_nvcmen_buf),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven_buf),
     .bgr(bgr), .bgr_int(bgr_int), .ngate_25(ngate_25),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv), .vpp(vpp),
     .vpp_int(vpp_int), .vpxa(vpxa), .vpxa_int(vpxa),
     .ysup_25(ysup_25), .vblinhi(vblinhi),
     .tm_testdec(fsm_tm_testdec));

endmodule
// Library - misc, Cell - nvcm_top, View - schematic
// LAST TIME SAVED: Feb 23 14:03:16 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module nvcm_top ( bp0, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_redrow,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_recall,
     fsm_rowadd, fsm_sample, fsm_tm_allbank_sel, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_dma,
     fsm_tm_margin0_read, fsm_tm_rd_mode, fsm_tm_tcol, fsm_tm_testdec,
     fsm_tm_testdec_wr, fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvpp, fsm_tm_xvpxa, fsm_tm_xvpxa_int,
     fsm_trim_ipp, fsm_trim_multibl_read, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_trim_vbg, fsm_trim_vpgmwl, fsm_trim_vrdwl,
     fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     nvcm_boot, nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b, clk,
     nv_dataout, nvcm_ce_b, nvcm_max_coladd, nvcm_max_rowadd, rst_b,
     smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_redrow, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_recall, fsm_sample, fsm_tm_allbank_sel,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_dma, fsm_tm_margin0_read, fsm_tm_rd_mode, fsm_tm_tcol,
     fsm_tm_testdec, fsm_tm_testdec_wr, fsm_tm_trow, fsm_tm_vwleqbl,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvpp, fsm_tm_xvpxa,
     fsm_tm_xvpxa_int, fsm_trim_multibl_read, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

output [11:0]  fsm_coladd;
output [2:0]  fsm_trim_vrdwl;
output [3:0]  fsm_blkadd;
output [2:0]  fsm_trim_rrefpgm;
output [3:0]  fsm_blkadd_b;
output [8:0]  fsm_rowadd;
output [2:0]  fsm_trim_rrefrd;
output [3:0]  fsm_trim_ipp;
output [3:0]  fsm_trim_vbg;
output [2:0]  fsm_trim_vpgmwl;

input [8:0]  nv_dataout;
input [8:0]  nvcm_max_rowadd;
input [11:0]  nvcm_max_coladd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - misc, Cell - nvcm_ml_block_1f, View - schematic
// LAST TIME SAVED: Feb 26 17:15:49 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module nvcm_ml_block_1f ( bp0, fsm_recall, fsm_tm_margin0_read,
     nvcm_boot, nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b, vpp,
     clk, nvcm_ce_b, nvcm_max_coladd, nvcm_max_rowadd, rst_b,
     smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_recall, fsm_tm_margin0_read, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b;

inout  vpp;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

input [11:0]  nvcm_max_coladd;
input [8:0]  nvcm_max_rowadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [8:0]  nv_dataout;

wire  [2:0]  fsm_trim_rrefpgm;

wire  [2:0]  fsm_trim_vrdwl;

wire  [11:0]  fsm_coladd;

wire  [3:0]  fsm_blkadd;

wire  [2:0]  fsm_trim_vpgmwl;

wire  [3:0]  fsm_trim_ipp;

wire  [2:0]  fsm_trim_rrefrd;

wire  [3:0]  fsm_blkadd_b;

wire  [3:0]  fsm_trim_vbg;

wire  [8:0]  fsm_rowadd;


/*
ml_chip_nvcm_1f Iml_chip_nvcm ( .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_coladd(fsm_coladd[8:0]), .tm_wleqbl(fsm_tm_vwleqbl),
     .tm_testdec_wr(fsm_tm_testdec_wr), .tm_tcol(fsm_tm_tcol),
     .tm_dma(fsm_tm_dma), .tm_allwl_l(fsm_tm_allwl_l),
     .tm_allwl_h(fsm_tm_allwl_h), .tm_allbl_l(fsm_tm_allbl_l),
     .tm_allbl_h(fsm_tm_allbl_h), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wren(fsm_wren), .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vrdwl(fsm_trim_vrdwl[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_vpgmwl(fsm_trim_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_xvpxaint(fsm_tm_xvpxa_int), .fsm_tm_xvpxa(fsm_tm_xvpxa),
     .fsm_tm_xvppint(fsm_tm_xvpp), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(rst_bd), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rrow(fsm_nv_redrow), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream),
     .fsm_multibl_read(fsm_trim_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_din(fsm_din),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .nv_dataout(nv_dataout[8:0]), .vpp(vpp));
sg_bufx10 I217 ( .in(rst_b), .out(rst_bd));
nvcm_top Invcm_top ( .fsm_coladd(fsm_coladd[11:0]),
     .nvcm_max_coladd(nvcm_max_coladd[11:0]),
     .nvcm_max_rowadd(nvcm_max_rowadd[8:0]),
     .fsm_tm_allbank_sel(fsm_tm_allbank_sel), .nvcm_boot(nvcm_boot),
     .spi_ss_b(spi_ss_b), .spi_sdi(spi_sdi),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .nvcm_ce_b(nvcm_ce_b), .nv_dataout(nv_dataout[8:0]), .clk(clk),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .nvcm_relextspi(nvcm_relextspi), .nvcm_rdy(nvcm_rdy),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_trim_vrdwl(fsm_trim_vrdwl[2:0]),
     .fsm_trim_vpgmwl(fsm_trim_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_multibl_read(fsm_trim_multibl_read),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_xvpxa_int(fsm_tm_xvpxa_int), .fsm_tm_xvpxa(fsm_tm_xvpxa),
     .fsm_tm_xvpp(fsm_tm_xvpp), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_vwleqbl(fsm_tm_vwleqbl), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_testdec_wr(fsm_tm_testdec_wr),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_tcol(fsm_tm_tcol),
     .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_margin0_read(fsm_tm_margin0_read),
     .fsm_tm_dma(fsm_tm_dma), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_sample(fsm_sample),
     .fsm_rowadd(fsm_rowadd[8:0]), .fsm_recall(fsm_recall),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_redrow(fsm_nv_redrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_din(fsm_din),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .bp0(bp0));
*/
endmodule
// Library - chip, Cell - nvcm_smc_fsm, View - schematic
// LAST TIME SAVED: May 29 16:32:39 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module nvcm_smc_fsm ( bm_banksel_i, bm_init_i, bm_rcapmux_en_i,
     bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bs_en0, cdone_out, ceb0, cm_banksel_blbrd_2_,
     cm_banksel_bldld, cm_banksel_bltrd_3_, cm_clk_blbrd, cm_sdi_u1,
     cm_sdi_u2d, cm_sdi_u3d, core_por_b0, core_por_bb, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_sdi_u0, cram_vddoff,
     cram_wl_en, cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b, end_of_startup, gint_hz, gsr, hiz_b0, j_rst_b,
     j_tck, j_tdi, md_spi_b, mode0, psdo, row_test0, sdo_enable,
     shift0, smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out_b, totdopad,
     update0, bm_sdo_o, cdone_in, cm_sdo_u0d1, cm_sdo_u1d3,
     cm_sdo_u2d1, cm_sdo_u3dd, creset_b_int, fabric_out_12_00,
     fabric_out_13_01, fabric_out_13_02, fromsdo, last_rsr3,
     monitor_celld4, .monitor_celldd(monitor_celld),
     smc_core_por_bottom1, smc_core_por_bottom2, spi_ss_in_bbankd,
     spi_ss_in_r, tck_pad, tdi_pad, tiegnd, tievdd, tms_pad, trst_pad,
     vpp );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, cm_banksel_bltrd_3_, cm_clk_blbrd,
     core_por_b0, core_por_bb, cram_pgateoff, cram_prec, cram_pullup_b,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, data_muxsel1_blbrd,
     data_muxsel_blbrd, en_8bconfig_b, end_of_startup, gint_hz, gsr,
     hiz_b0, j_rst_b, j_tck, j_tdi, md_spi_b, mode0, row_test0,
     sdo_enable, shift0, smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd,
     smc_write, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out_b,
     totdopad, update0;

input  cdone_in, creset_b_int, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fromsdo, last_rsr3, smc_core_por_bottom1,
     smc_core_por_bottom2, tck_pad, tdi_pad, tiegnd, tievdd, tms_pad,
     trst_pad, vpp;

output [7:0]  bm_sa_i;
output [1:0]  cram_sdi_u0;
output [1:0]  cm_sdi_u2d;
output [1:0]  cm_banksel_bldld;
output [3:0]  bm_banksel_i;
output [1:0]  cm_sdi_u1;
output [1:0]  cm_sdi_u3d;
output [7:1]  psdo;
output [3:0]  bm_sdi_i;

input [3:2]  monitor_celld;
input [7:1]  spi_ss_in_r;
input [1:0]  cm_sdo_u0d1;
input [3:0]  bm_sdo_o;
input [1:0]  cm_sdo_u3dd;
input [1:0]  cm_sdo_u1d3;
input [1:0]  cm_sdo_u2d1;
input [4:0]  spi_ss_in_bbankd;
input [1:0]  monitor_celld4;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  cm_banksel_nbuf;



CHIP_smc_ice12k Ismc_ice1f ( .vddio_rightbank(vddp_),
     .trst_pad(trst_pad), .tms_pad(tms_pad), .tdi_pad(tdi_pad),
     .tck_pad(tck_pad), .spi_ss_in_r(spi_ss_in_r[7:1]),
     .spi_ss_in_bbank(spi_ss_in_bbankd[4:0]),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_spi_sdo(nvcm_spi_sdo), .nvcm_relextspi(nvcm_relextspi),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot),
     .monitor_celld(monitor_celld[3:2]),
     .monitor_celld4(monitor_celld4[1:0]), .last_rsr3(last_rsr3),
     .idcode_msb20bits({tiegnd, tiegnd, tiegnd, tievdd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tievdd}),
     .fromsdo(fromsdo), .fabric_out_41_02(fabric_out_13_02),
     .fabric_out_41_01(fabric_out_13_01),
     .fabric_out_40_00(fabric_out_12_00),
     .cm_sdo_u3d1(cm_sdo_u3dd[1:0]), .cm_sdo_u2d1(cm_sdo_u2d1[1:0]),
     .cm_sdo_u1d3(cm_sdo_u1d3[1:0]), .cm_sdo_u0d1(cm_sdo_u0d1[1:0]),
     .cdone_in(cdone_in), .bp0(bp0), .bm_sdo_o(bm_sdo_o[3:0]),
     .update0(update0), .totdopad(totdopad),
     .spi_ss_out_b(spi_ss_out_b), .spi_sdo_oe_b(spi_sdo_oe_b),
     .spi_sdo(spi_sdo), .spi_clk_out(spi_clk_out),
     .smc_write0(smc_write), .smc_wdis_dclk(smc_wdis_dclk_blbrd),
     .smc_rsr_rst(smc_rsr_rst), .smc_row_inc(smc_row_inc),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream),
     .smc_clk_out(cm_clk_blbrd), .shift0(shift0),
     .sdo_enable(sdo_enable), .rst_b(rst_b_4smc2nvcm),
     .row_test0(row_test0), .psdo(psdo[7:1]),
     .nvcm_spi_ss_b(nvcm_spi_ss_b), .nvcm_spi_sdi(nvcm_spi_sdi),
     .mode0(mode0), .md_spi_b(md_spi_b), .j_tdi(j_tdi), .j_tck(j_tck),
     .j_rst_b(j_rst_b), .hiz_b0(hiz_b0), .gsr(gsr), .gint_hz(gint_hz),
     .end_of_startup(end_of_startup), .en_8bconfig_b(en_8bconfig_b),
     .data_muxsel1(data_muxsel1_blbrd),
     .data_muxsel(data_muxsel_blbrd), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_pgateoff(cram_pgateoff),
     .core_por_bb(core_por_bb), .core_por_b0(core_por_b0),
     .cm_sdi_u3(cm_sdi_u3d[1:0]), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u0(cram_sdi_u0[1:0]),
     .cm_banksel_bldld(cm_banksel_bldld[1:0]),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_),
     .cm_banksel({cm_banksel_bltrd_3_, cm_banksel_nbuf[2:0]}),
     .ceb0(ceb0), .cdone_out(cdone_out), .bs_en0(bs_en0),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .bm_banksel_i(bm_banksel_i[3:0]),
     .creset_b_int(creset_b_int));
nvcm_ml_block_1f Invcm_ml_block_1f ( .nvcm_max_coladd({tiegnd, tiegnd,
     tiegnd, tievdd, tiegnd, tievdd, tiegnd, tiegnd, tiegnd, tievdd,
     tievdd, tievdd}), .nvcm_max_rowadd({tiegnd, tiegnd, tievdd,
     tievdd, tiegnd, tiegnd, tievdd, tievdd, tievdd}),
     .spi_ss_b(nvcm_spi_ss_b), .spi_sdi(nvcm_spi_sdi),
     .rst_b(rst_b_4smc2nvcm), .nvcm_ce_b(end_of_startup),
     .clk(spi_clk_out), .spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .spi_sdo(nvcm_spi_sdo), .nvcm_rdy(nvcm_rdy),
     .nvcm_boot(nvcm_boot),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream),
     .fsm_tm_margin0_read(net260), .fsm_recall(net261), .bp0(bp0),
     .nvcm_relextspi(nvcm_relextspi), .vpp(vpp));

endmodule
// Library - xpmem, Cell - ml_buf_ice5_2, View - schematic
// LAST TIME SAVED: Aug 15 18:07:29 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_buf_ice5_2 ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));
inv_hvt I391 ( .A(net77), .Y(o));

endmodule
// Library - io, Cell - topbank_1k_july16, View - schematic
// LAST TIME SAVED: Jul 21 09:24:34 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module topbank_1k_july16 ( in, pad, vpp, vppin, oen, out, ren );

inout  vpp, vppin;


output [23:0]  in;

inout [23:0]  pad;

input [23:0]  oen;
input [23:0]  ren;
input [23:0]  out;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



PVDD2POC I66 ( .VDDPST(vddio_topbank));
pvpp I62 ( .vppin(vppin), .vpp(vpp));
PDUW08DGZ I46_9_ ( .PAD(pad[9]), .C(in[9]), .OEN(oen[9]), .I(out[9]),
     .REN(ren[9]));
PDUW08DGZ I46_8_ ( .PAD(pad[8]), .C(in[8]), .OEN(oen[8]), .I(out[8]),
     .REN(ren[8]));
PDUW08DGZ I46_7_ ( .PAD(pad[7]), .C(in[7]), .OEN(oen[7]), .I(out[7]),
     .REN(ren[7]));
PDUW08DGZ I46_6_ ( .PAD(pad[6]), .C(in[6]), .OEN(oen[6]), .I(out[6]),
     .REN(ren[6]));
PDUW08DGZ I46_5_ ( .PAD(pad[5]), .C(in[5]), .OEN(oen[5]), .I(out[5]),
     .REN(ren[5]));
PDUW08DGZ I46_4_ ( .PAD(pad[4]), .C(in[4]), .OEN(oen[4]), .I(out[4]),
     .REN(ren[4]));
PDUW08DGZ I50_12_ ( .PAD(pad[12]), .C(in[12]), .OEN(oen[12]),
     .I(out[12]), .REN(ren[12]));
PDUW08DGZ I50_11_ ( .PAD(pad[11]), .C(in[11]), .OEN(oen[11]),
     .I(out[11]), .REN(ren[11]));
PDUW08DGZ I73_10_ ( .PAD(pad[10]), .C(in[10]), .OEN(oen[10]),
     .I(out[10]), .REN(ren[10]));
PDUW08DGZ I71_16_ ( .PAD(pad[16]), .C(in[16]), .OEN(oen[16]),
     .I(out[16]), .REN(ren[16]));
PDUW08DGZ I71_15_ ( .PAD(pad[15]), .C(in[15]), .OEN(oen[15]),
     .I(out[15]), .REN(ren[15]));
PDUW08DGZ I71_14_ ( .PAD(pad[14]), .C(in[14]), .OEN(oen[14]),
     .I(out[14]), .REN(ren[14]));
PDUW08DGZ I71_13_ ( .PAD(pad[13]), .C(in[13]), .OEN(oen[13]),
     .I(out[13]), .REN(ren[13]));
PDUW08DGZ I51_23_ ( .PAD(pad[23]), .C(in[23]), .OEN(oen[23]),
     .I(out[23]), .REN(ren[23]));
PDUW08DGZ I51_22_ ( .PAD(pad[22]), .C(in[22]), .OEN(oen[22]),
     .I(out[22]), .REN(ren[22]));
PDUW08DGZ I51_21_ ( .PAD(pad[21]), .C(in[21]), .OEN(oen[21]),
     .I(out[21]), .REN(ren[21]));
PDUW08DGZ I51_20_ ( .PAD(pad[20]), .C(in[20]), .OEN(oen[20]),
     .I(out[20]), .REN(ren[20]));
PDUW08DGZ I51_19_ ( .PAD(pad[19]), .C(in[19]), .OEN(oen[19]),
     .I(out[19]), .REN(ren[19]));
PDUW08DGZ I51_18_ ( .PAD(pad[18]), .C(in[18]), .OEN(oen[18]),
     .I(out[18]), .REN(ren[18]));
PDUW08DGZ I51_17_ ( .PAD(pad[17]), .C(in[17]), .OEN(oen[17]),
     .I(out[17]), .REN(ren[17]));
PDUW08DGZ I42_3_ ( .PAD(pad[3]), .C(in[3]), .OEN(oen[3]), .I(out[3]),
     .REN(ren[3]));
PDUW08DGZ I42_2_ ( .PAD(pad[2]), .C(in[2]), .OEN(oen[2]), .I(out[2]),
     .REN(ren[2]));
PDUW08DGZ I42_1_ ( .PAD(pad[1]), .C(in[1]), .OEN(oen[1]), .I(out[1]),
     .REN(ren[1]));
PDUW08DGZ I42_0_ ( .PAD(pad[0]), .C(in[0]), .OEN(oen[0]), .I(out[0]),
     .REN(ren[0]));
PVDD1DGZ I58_1_ ( .VDD(vdd_));
PVDD1DGZ I58_0_ ( .VDD(vdd_));
PVDD2DGZ I57_1_ ( .VDDPST(vddio_topbank));
PVDD2DGZ I57_0_ ( .VDDPST(vddio_topbank));
PVDD2DGZ I72_1_ ( .VDDPST(vddio_topbank));
PVDD2DGZ I72_0_ ( .VDDPST(vddio_topbank));
PVSS3DGZ I32 ( .VSS(gnd_));
PVSS3DGZ I70_1_ ( .VSS(gnd_));
PVSS3DGZ I70_0_ ( .VSS(gnd_));
PVSS3DGZ I68_1_ ( .VSS(gnd_));
PVSS3DGZ I68_0_ ( .VSS(gnd_));

endmodule
// Library - xpmem, Cell - ml_rowdrv2_last, View - schematic
// LAST TIME SAVED: Sep 26 14:07:07 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_rowdrv2_last ( pgate, reset, smc_rsr_out, vddctrl, wl,
     wl_rd_sup, wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write
     );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  NM0 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
ml_dff_schematic I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));

endmodule
// Library - xpmem, Cell - ml_rowdrvsup2, View - schematic
// LAST TIME SAVED: Oct  6 17:48:55 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_rowdrvsup2 ( wl_rd_sup, wl_rden_b );
inout  wl_rd_sup, wl_rden_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



tielo I228 ( .tielo(net0140));
rppolywo_m  R10 ( .MINUS(net045), .PLUS(net0110), .BULK(gnd_));
rppolywo_m  R14 ( .MINUS(wl_rd_sup), .PLUS(net0113), .BULK(gnd_));
rppolywo_m  R12 ( .MINUS(net0104), .PLUS(wl_rd_sup), .BULK(gnd_));
rppolywo_m  R13 ( .MINUS(net0107), .PLUS(net0108), .BULK(gnd_));
rppolywo_m  R11 ( .MINUS(net0110), .PLUS(net0104), .BULK(gnd_));
rppolywo_m  R15 ( .MINUS(net0113), .PLUS(net0107), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(net071), .PLUS(net077), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net0108), .PLUS(net071), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(net077), .PLUS(net083), .BULK(gnd_));
rppolywo_m  R19 ( .MINUS(net080), .PLUS(net092), .BULK(gnd_));
rppolywo_m  R20 ( .MINUS(net083), .PLUS(net086), .BULK(gnd_));
rppolywo_m  R21 ( .MINUS(net086), .PLUS(net080), .BULK(gnd_));
rppolywo_m  R22 ( .MINUS(net089), .PLUS(net095), .BULK(gnd_));
rppolywo_m  R23 ( .MINUS(net092), .PLUS(net089), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(net095), .PLUS(net0158), .BULK(gnd_));
inv_hvt I217 ( .A(wl_rden_b), .Y(net0142));
inv_hvt I220 ( .A(net0142), .Y(act_rd_b));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
nch_hvt  MN16 ( .D(wl_rd_sup), .B(gnd_), .G(act_rd_b), .S(gnd_));
nch_hvt  MN14 ( .D(net0158), .B(gnd_), .G(act_rd), .S(gnd_));
pch_hvt  MP13 ( .D(wl_rden_b), .B(vdd_), .G(net0140), .S(vdd_));
pch_hvt  MP15 ( .D(net045), .B(vdd_), .G(act_rd_b), .S(vdd_));

endmodule
// Library - xpmem, Cell - ml_rowdrv2, View - schematic
// LAST TIME SAVED: Aug 23 15:16:05 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_rowdrv2 ( pgate, reset, smc_rsr_out, vddctrl, wl, wl_rd_sup,
     wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
ml_dff_schematic I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile_last, View - schematic
// LAST TIME SAVED: Aug  9 15:08:40 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_rowdrv_tile_last ( pgate, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  wl;
output [15:0]  reset;
output [15:0]  pgate;
output [15:0]  vddctrl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  smc_rsr_out;



nor2_hvt I211 ( .A(smc_rsr_out[15]), .Y(net049), .B(smc_rsr_inc_out));
ml_rowdrv2_last Iml_rowdrv2_last ( .smc_rsr_inc(smc_rsr_inc_last),
     .smc_rsr_in(smc_rsr_out[14]), .rsr_rst(rsr_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_rst(cram_rst_buf),
     .smc_rsr_out(smc_rsr_out[15]), .reset(reset[15]), .wl(wl[15]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]));
inv_hvt I391 ( .A(net049), .Y(smc_rsr_inc_last));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I194 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I195 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I198 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I207 ( .A(net041), .Y(por_rst_buf));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net079));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I200 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I206 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I190 ( .A(net079), .Y(smc_rsr_1st_out));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile, View - schematic
// LAST TIME SAVED: Aug 15 11:21:19 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_rowdrv_tile ( pgate, por_rst_out, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  por_rst_out, smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  vddctrl;
output [15:0]  reset;
output [15:0]  pgate;
output [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  smc_rsr_out;



inv_hvt I207 ( .A(net041), .Y(por_rst_out));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I194 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I195 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I198 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I190 ( .A(net037), .Y(smc_rsr_1st_out));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net037));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I200 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I206 ( .A(net047), .Y(rsr_rst_buf));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_15_ ( .reset(reset[15]), .wl(wl[15]),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[14]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[15]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_rowdrv_bank_1k, View - schematic
// LAST TIME SAVED: Mar  9 16:48:31 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_rowdrv_bank_1k ( jtag_rowtest_mode_b, last_rsr, pgate, reset,
     vddctrl, wl, banksel, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst,
     smc_rsr_inc, smc_write, trst_b );
output  jtag_rowtest_mode_b, last_rsr;

input  banksel, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst, smc_rsr_inc,
     smc_write, trst_b;

output [143:0]  reset;
output [143:0]  wl;
output [143:0]  pgate;
output [143:0]  vddctrl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  smc_rsr_1st_out_buf;

wire  [8:0]  smc_rsr_out;

wire  [7:0]  por_rst_out;

wire  [7:0]  smc_rsr_inc_out;

wire  [0:8]  smc_rsr_1st_out;



vdd_tielow I251 ( .gnd_tiel(net0130));
tiehi I269 ( .tiehi(net162));
tiehi I249 ( .tiehi(net131));
tiehi I250 ( .tiehi(net132));
ml_buf_ice5_2 I227 ( .in(net131), .o(net134), .sel(net131));
ml_buf_ice5_2 I216 ( .in(net131), .o(net137), .sel(net131));
ml_buf_ice5_2 I198 ( .sel(banksel), .in(cram_wl_en),
     .o(cram_wl_en_buf));
ml_buf_ice5_2 I196 ( .sel(banksel), .in(cram_rst), .o(cram_rst_buf));
ml_buf_ice5_2 I199 ( .sel(net132), .in(por_rst), .o(por_rst_buf));
ml_buf_ice5_2 I197 ( .sel(banksel), .in(cram_vddoff),
     .o(cram_vddoff_buf));
ml_buf_ice5_2 I195 ( .sel(banksel), .in(cram_pgateoff),
     .o(cram_pgateoff_buf));
ml_buf_ice5_2 I201 ( .sel(banksel), .in(smc_write), .o(smc_write_buf));
ml_buf_ice5_2 I203 ( .sel(net184), .in(net184), .o(smc_rsr_inc_buf));
ml_buf_ice5_2 I213 ( .in(net162), .o(net161), .sel(net162));
ml_rowdrv_tile_last Iml_rowdrv_tile_last (
     .smc_rsr_inc_out(smc_rsr_inc_out_last), .pgate(pgate[143:128]),
     .wl(wl[143:128]), .vddctrl(vddctrl[143:128]),
     .reset(reset[143:128]), .smc_rsr_1st_out(smc_rsr_1st_out[8]),
     .smcc_rsr_out(smc_rsr_out[8]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_buf), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[7]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf));
nand2_hvt I233 ( .A(smc_rsr_inc), .B(banksel), .Y(net181));
mux2_hvt I161 ( .in1(jtag_clk), .in0(net263), .out(net184),
     .sel(net256));
nand3_hvt I231 ( .Y(net186), .B(net190), .C(net190), .A(net190));
nand3_hvt I230 ( .Y(net190), .B(net195), .C(net195), .A(net195));
nand3_hvt I224 ( .B(net131), .Y(net195), .A(net131), .C(net131));
nor3_hvt I238 ( .B(por_rst), .Y(net248), .A(net208), .C(trst));
nor3_hvt I232 ( .C(rsr_rst), .A(jtag_rowtest_rst), .B(net0130),
     .Y(net213));
nor3_hvt I218 ( .B(net225), .Y(net215), .A(net225), .C(net225));
nor3_hvt I220 ( .B(net215), .Y(net219), .A(net215), .C(net215));
nor3_hvt I217 ( .C(net131), .A(net131), .B(net131), .Y(net225));
nor3_hvt I244 ( .B(por_rst), .Y(net227), .A(net276),
     .C(smc_rsr_1st_out_buf[0]));
ml_rowdrv_tile Iml_rowdrv_tile_7_ ( .por_rst_out(por_rst_out[7]),
     .smc_rsr_inc_out(smc_rsr_inc_out[7]),
     .smcc_rsr_out(smc_rsr_out[7]),
     .smc_rsr_1st_out(smc_rsr_1st_out[7]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out_last), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[6]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[127:112]), .vddctrl(vddctrl[127:112]),
     .reset(reset[127:112]), .pgate(pgate[127:112]));
ml_rowdrv_tile Iml_rowdrv_tile_6_ ( .por_rst_out(por_rst_out[6]),
     .smc_rsr_inc_out(smc_rsr_inc_out[6]),
     .smcc_rsr_out(smc_rsr_out[6]),
     .smc_rsr_1st_out(smc_rsr_1st_out[6]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[7]), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[5]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[111:96]), .vddctrl(vddctrl[111:96]), .reset(reset[111:96]),
     .pgate(pgate[111:96]));
ml_rowdrv_tile Iml_rowdrv_tile_5_ ( .por_rst_out(por_rst_out[5]),
     .smc_rsr_inc_out(smc_rsr_inc_out[5]),
     .smcc_rsr_out(smc_rsr_out[5]),
     .smc_rsr_1st_out(smc_rsr_1st_out[5]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[6]), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[4]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[95:80]), .vddctrl(vddctrl[95:80]), .reset(reset[95:80]),
     .pgate(pgate[95:80]));
ml_rowdrv_tile Iml_rowdrv_tile_4_ ( .por_rst_out(por_rst_out[4]),
     .smc_rsr_inc_out(smc_rsr_inc_out[4]),
     .smcc_rsr_out(smc_rsr_out[4]),
     .smc_rsr_1st_out(smc_rsr_1st_out[4]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[5]), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[3]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[79:64]), .vddctrl(vddctrl[79:64]), .reset(reset[79:64]),
     .pgate(pgate[79:64]));
ml_rowdrv_tile Iml_rowdrv_tile_3_ ( .por_rst_out(por_rst_out[3]),
     .smc_rsr_inc_out(smc_rsr_inc_out[3]),
     .smcc_rsr_out(smc_rsr_out[3]),
     .smc_rsr_1st_out(smc_rsr_1st_out[3]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[4]), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[2]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[63:48]), .vddctrl(vddctrl[63:48]), .reset(reset[63:48]),
     .pgate(pgate[63:48]));
ml_rowdrv_tile Iml_rowdrv_tile_2_ ( .por_rst_out(por_rst_out[2]),
     .smc_rsr_inc_out(smc_rsr_inc_out[2]),
     .smcc_rsr_out(smc_rsr_out[2]),
     .smc_rsr_1st_out(smc_rsr_1st_out[2]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[3]), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[1]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[47:32]), .vddctrl(vddctrl[47:32]), .reset(reset[47:32]),
     .pgate(pgate[47:32]));
ml_rowdrv_tile Iml_rowdrv_tile_1_ ( .por_rst_out(por_rst_out[1]),
     .smc_rsr_inc_out(smc_rsr_inc_out[1]),
     .smcc_rsr_out(smc_rsr_out[1]),
     .smc_rsr_1st_out(smc_rsr_1st_out[1]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[2]), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[0]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[31:16]), .vddctrl(vddctrl[31:16]), .reset(reset[31:16]),
     .pgate(pgate[31:16]));
ml_rowdrv_tile Iml_rowdrv_tile_0_ ( .por_rst_out(por_rst_out[0]),
     .smc_rsr_inc_out(smc_rsr_inc_out[0]),
     .smcc_rsr_out(smc_rsr_out[0]),
     .smc_rsr_1st_out(smc_rsr_1st_out[0]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[1]), .smc_rsr_in(smc_rsr_in_1st),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[15:0]), .vddctrl(vddctrl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]));
nor2_hvt I239 ( .A(jtag_rowtest_rst), .B(net248), .Y(net208));
nor2_hvt I193 ( .A(por_rst), .B(rsr_set_1st), .Y(net252));
nor2_hvt I245 ( .A(rsr_set_1st), .B(net227), .Y(net276));
inv_hvt I247 ( .A(net256), .Y(jtag_rowtest_mode_b));
inv_hvt I241 ( .A(net208), .Y(net256));
inv_hvt I192 ( .A(net213), .Y(rsr_set_1st));
inv_hvt I234 ( .A(net181), .Y(net263));
inv_hvt I35 ( .A(net264), .Y(smc_rsr_1st_out_buf[0]));
inv_hvt I240 ( .A(trst_b), .Y(trst));
inv_hvt I210 ( .A(net268), .Y(last_rsr));
inv_hvt I391 ( .A(net252), .Y(rst_row_reg));
inv_hvt I36 ( .A(smc_rsr_1st_out[0]), .Y(net264));
inv_hvt I209 ( .A(smc_rsr_out[8]), .Y(net268));
inv_hvt I205 ( .A(net276), .Y(smc_rsr_in_1st));

endmodule
// Library - leafcell, Cell - bram_bufferx4, View - schematic
// LAST TIME SAVED: Jun 25 13:46:30 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module bram_bufferx4 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - xpmem, Cell - sg_dffbuf_modified, View - schematic
// LAST TIME SAVED: Jun 12 15:50:42 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module sg_dffbuf_modified ( dffout, clk, d, r );
output  dffout;

input  clk, d, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I2 ( .in(net10), .out(dffout));
ml_dff I0 ( .R(r), .D(d), .CLK(clk), .QN(net9), .Q(net10));

endmodule
// Library - chip, Cell - CHIP_route_left1f, View - schematic
// LAST TIME SAVED: May 12 08:56:33 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module CHIP_route_left1f ( cm_banksel_bltld3_1_, cm_clk_bltld3,
     cm_sdi_u1d3[1:0], cm_sdo_u1d1[1:0], core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, last_rsr[1:0],
     monitor_celld2[1:0], pgate_l[287:0], reset_l[287:0],
     smc_wdis_dclk_bltld3, vdd_cntl_l[287:0], wl_l[287:0],
     cf_lbank[300], cf_lbank[479], cm_banksel_blbld1[0],
     cm_banksel_blbld[1], cm_clk_blbld, cm_sdi_u1d[1:0],
     cm_sdo_u1[1:0], core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0 );
output  cm_banksel_bltld3_1_, cm_clk_bltld3, core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, smc_wdis_dclk_bltld3;

input  cm_clk_blbld, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;

output [1:0]  last_rsr;
output [1:0]  cm_sdo_u1d1;
output [1:0]  cm_sdi_u1d3;
output [287:0]  reset_l;
output [1:0]  monitor_celld2;
output [287:0]  vdd_cntl_l;
output [287:0]  pgate_l;
output [287:0]  wl_l;

input [1:0]  cm_sdi_u1d;
input [300:479]  cf_lbank;
input [1:1]  cm_banksel_blbld;
input [1:0]  cm_sdo_u1;
input [0:0]  cm_banksel_blbld1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u1d0;

wire  [1:0]  cm_sdo_u1d;

wire  [1:0]  cm_sdi_u1d0;

wire  [0:1]  net129;

wire  [1:0]  dff_out;

wire  [1:1]  monitor_celld1;

wire  [1:1]  monitor_celld;

wire  [1:1]  cm_banksel_bltld;



ml_rowdrv_bank_1k Irowul ( .vddctrl({vdd_cntl_l[144], vdd_cntl_l[145],
     vdd_cntl_l[146], vdd_cntl_l[147], vdd_cntl_l[148],
     vdd_cntl_l[149], vdd_cntl_l[150], vdd_cntl_l[151],
     vdd_cntl_l[152], vdd_cntl_l[153], vdd_cntl_l[154],
     vdd_cntl_l[155], vdd_cntl_l[156], vdd_cntl_l[157],
     vdd_cntl_l[158], vdd_cntl_l[159], vdd_cntl_l[160],
     vdd_cntl_l[161], vdd_cntl_l[162], vdd_cntl_l[163],
     vdd_cntl_l[164], vdd_cntl_l[165], vdd_cntl_l[166],
     vdd_cntl_l[167], vdd_cntl_l[168], vdd_cntl_l[169],
     vdd_cntl_l[170], vdd_cntl_l[171], vdd_cntl_l[172],
     vdd_cntl_l[173], vdd_cntl_l[174], vdd_cntl_l[175],
     vdd_cntl_l[176], vdd_cntl_l[177], vdd_cntl_l[178],
     vdd_cntl_l[179], vdd_cntl_l[180], vdd_cntl_l[181],
     vdd_cntl_l[182], vdd_cntl_l[183], vdd_cntl_l[184],
     vdd_cntl_l[185], vdd_cntl_l[186], vdd_cntl_l[187],
     vdd_cntl_l[188], vdd_cntl_l[189], vdd_cntl_l[190],
     vdd_cntl_l[191], vdd_cntl_l[192], vdd_cntl_l[193],
     vdd_cntl_l[194], vdd_cntl_l[195], vdd_cntl_l[196],
     vdd_cntl_l[197], vdd_cntl_l[198], vdd_cntl_l[199],
     vdd_cntl_l[200], vdd_cntl_l[201], vdd_cntl_l[202],
     vdd_cntl_l[203], vdd_cntl_l[204], vdd_cntl_l[205],
     vdd_cntl_l[206], vdd_cntl_l[207], vdd_cntl_l[208],
     vdd_cntl_l[209], vdd_cntl_l[210], vdd_cntl_l[211],
     vdd_cntl_l[212], vdd_cntl_l[213], vdd_cntl_l[214],
     vdd_cntl_l[215], vdd_cntl_l[216], vdd_cntl_l[217],
     vdd_cntl_l[218], vdd_cntl_l[219], vdd_cntl_l[220],
     vdd_cntl_l[221], vdd_cntl_l[222], vdd_cntl_l[223],
     vdd_cntl_l[224], vdd_cntl_l[225], vdd_cntl_l[226],
     vdd_cntl_l[227], vdd_cntl_l[228], vdd_cntl_l[229],
     vdd_cntl_l[230], vdd_cntl_l[231], vdd_cntl_l[232],
     vdd_cntl_l[233], vdd_cntl_l[234], vdd_cntl_l[235],
     vdd_cntl_l[236], vdd_cntl_l[237], vdd_cntl_l[238],
     vdd_cntl_l[239], vdd_cntl_l[240], vdd_cntl_l[241],
     vdd_cntl_l[242], vdd_cntl_l[243], vdd_cntl_l[244],
     vdd_cntl_l[245], vdd_cntl_l[246], vdd_cntl_l[247],
     vdd_cntl_l[248], vdd_cntl_l[249], vdd_cntl_l[250],
     vdd_cntl_l[251], vdd_cntl_l[252], vdd_cntl_l[253],
     vdd_cntl_l[254], vdd_cntl_l[255], vdd_cntl_l[256],
     vdd_cntl_l[257], vdd_cntl_l[258], vdd_cntl_l[259],
     vdd_cntl_l[260], vdd_cntl_l[261], vdd_cntl_l[262],
     vdd_cntl_l[263], vdd_cntl_l[264], vdd_cntl_l[265],
     vdd_cntl_l[266], vdd_cntl_l[267], vdd_cntl_l[268],
     vdd_cntl_l[269], vdd_cntl_l[270], vdd_cntl_l[271],
     vdd_cntl_l[272], vdd_cntl_l[273], vdd_cntl_l[274],
     vdd_cntl_l[275], vdd_cntl_l[276], vdd_cntl_l[277],
     vdd_cntl_l[278], vdd_cntl_l[279], vdd_cntl_l[280],
     vdd_cntl_l[281], vdd_cntl_l[282], vdd_cntl_l[283],
     vdd_cntl_l[284], vdd_cntl_l[285], vdd_cntl_l[286],
     vdd_cntl_l[287]}), .wl({wl_l[144], wl_l[145], wl_l[146],
     wl_l[147], wl_l[148], wl_l[149], wl_l[150], wl_l[151], wl_l[152],
     wl_l[153], wl_l[154], wl_l[155], wl_l[156], wl_l[157], wl_l[158],
     wl_l[159], wl_l[160], wl_l[161], wl_l[162], wl_l[163], wl_l[164],
     wl_l[165], wl_l[166], wl_l[167], wl_l[168], wl_l[169], wl_l[170],
     wl_l[171], wl_l[172], wl_l[173], wl_l[174], wl_l[175], wl_l[176],
     wl_l[177], wl_l[178], wl_l[179], wl_l[180], wl_l[181], wl_l[182],
     wl_l[183], wl_l[184], wl_l[185], wl_l[186], wl_l[187], wl_l[188],
     wl_l[189], wl_l[190], wl_l[191], wl_l[192], wl_l[193], wl_l[194],
     wl_l[195], wl_l[196], wl_l[197], wl_l[198], wl_l[199], wl_l[200],
     wl_l[201], wl_l[202], wl_l[203], wl_l[204], wl_l[205], wl_l[206],
     wl_l[207], wl_l[208], wl_l[209], wl_l[210], wl_l[211], wl_l[212],
     wl_l[213], wl_l[214], wl_l[215], wl_l[216], wl_l[217], wl_l[218],
     wl_l[219], wl_l[220], wl_l[221], wl_l[222], wl_l[223], wl_l[224],
     wl_l[225], wl_l[226], wl_l[227], wl_l[228], wl_l[229], wl_l[230],
     wl_l[231], wl_l[232], wl_l[233], wl_l[234], wl_l[235], wl_l[236],
     wl_l[237], wl_l[238], wl_l[239], wl_l[240], wl_l[241], wl_l[242],
     wl_l[243], wl_l[244], wl_l[245], wl_l[246], wl_l[247], wl_l[248],
     wl_l[249], wl_l[250], wl_l[251], wl_l[252], wl_l[253], wl_l[254],
     wl_l[255], wl_l[256], wl_l[257], wl_l[258], wl_l[259], wl_l[260],
     wl_l[261], wl_l[262], wl_l[263], wl_l[264], wl_l[265], wl_l[266],
     wl_l[267], wl_l[268], wl_l[269], wl_l[270], wl_l[271], wl_l[272],
     wl_l[273], wl_l[274], wl_l[275], wl_l[276], wl_l[277], wl_l[278],
     wl_l[279], wl_l[280], wl_l[281], wl_l[282], wl_l[283], wl_l[284],
     wl_l[285], wl_l[286], wl_l[287]}), .reset({reset_l[144],
     reset_l[145], reset_l[146], reset_l[147], reset_l[148],
     reset_l[149], reset_l[150], reset_l[151], reset_l[152],
     reset_l[153], reset_l[154], reset_l[155], reset_l[156],
     reset_l[157], reset_l[158], reset_l[159], reset_l[160],
     reset_l[161], reset_l[162], reset_l[163], reset_l[164],
     reset_l[165], reset_l[166], reset_l[167], reset_l[168],
     reset_l[169], reset_l[170], reset_l[171], reset_l[172],
     reset_l[173], reset_l[174], reset_l[175], reset_l[176],
     reset_l[177], reset_l[178], reset_l[179], reset_l[180],
     reset_l[181], reset_l[182], reset_l[183], reset_l[184],
     reset_l[185], reset_l[186], reset_l[187], reset_l[188],
     reset_l[189], reset_l[190], reset_l[191], reset_l[192],
     reset_l[193], reset_l[194], reset_l[195], reset_l[196],
     reset_l[197], reset_l[198], reset_l[199], reset_l[200],
     reset_l[201], reset_l[202], reset_l[203], reset_l[204],
     reset_l[205], reset_l[206], reset_l[207], reset_l[208],
     reset_l[209], reset_l[210], reset_l[211], reset_l[212],
     reset_l[213], reset_l[214], reset_l[215], reset_l[216],
     reset_l[217], reset_l[218], reset_l[219], reset_l[220],
     reset_l[221], reset_l[222], reset_l[223], reset_l[224],
     reset_l[225], reset_l[226], reset_l[227], reset_l[228],
     reset_l[229], reset_l[230], reset_l[231], reset_l[232],
     reset_l[233], reset_l[234], reset_l[235], reset_l[236],
     reset_l[237], reset_l[238], reset_l[239], reset_l[240],
     reset_l[241], reset_l[242], reset_l[243], reset_l[244],
     reset_l[245], reset_l[246], reset_l[247], reset_l[248],
     reset_l[249], reset_l[250], reset_l[251], reset_l[252],
     reset_l[253], reset_l[254], reset_l[255], reset_l[256],
     reset_l[257], reset_l[258], reset_l[259], reset_l[260],
     reset_l[261], reset_l[262], reset_l[263], reset_l[264],
     reset_l[265], reset_l[266], reset_l[267], reset_l[268],
     reset_l[269], reset_l[270], reset_l[271], reset_l[272],
     reset_l[273], reset_l[274], reset_l[275], reset_l[276],
     reset_l[277], reset_l[278], reset_l[279], reset_l[280],
     reset_l[281], reset_l[282], reset_l[283], reset_l[284],
     reset_l[285], reset_l[286], reset_l[287]}), .pgate({pgate_l[144],
     pgate_l[145], pgate_l[146], pgate_l[147], pgate_l[148],
     pgate_l[149], pgate_l[150], pgate_l[151], pgate_l[152],
     pgate_l[153], pgate_l[154], pgate_l[155], pgate_l[156],
     pgate_l[157], pgate_l[158], pgate_l[159], pgate_l[160],
     pgate_l[161], pgate_l[162], pgate_l[163], pgate_l[164],
     pgate_l[165], pgate_l[166], pgate_l[167], pgate_l[168],
     pgate_l[169], pgate_l[170], pgate_l[171], pgate_l[172],
     pgate_l[173], pgate_l[174], pgate_l[175], pgate_l[176],
     pgate_l[177], pgate_l[178], pgate_l[179], pgate_l[180],
     pgate_l[181], pgate_l[182], pgate_l[183], pgate_l[184],
     pgate_l[185], pgate_l[186], pgate_l[187], pgate_l[188],
     pgate_l[189], pgate_l[190], pgate_l[191], pgate_l[192],
     pgate_l[193], pgate_l[194], pgate_l[195], pgate_l[196],
     pgate_l[197], pgate_l[198], pgate_l[199], pgate_l[200],
     pgate_l[201], pgate_l[202], pgate_l[203], pgate_l[204],
     pgate_l[205], pgate_l[206], pgate_l[207], pgate_l[208],
     pgate_l[209], pgate_l[210], pgate_l[211], pgate_l[212],
     pgate_l[213], pgate_l[214], pgate_l[215], pgate_l[216],
     pgate_l[217], pgate_l[218], pgate_l[219], pgate_l[220],
     pgate_l[221], pgate_l[222], pgate_l[223], pgate_l[224],
     pgate_l[225], pgate_l[226], pgate_l[227], pgate_l[228],
     pgate_l[229], pgate_l[230], pgate_l[231], pgate_l[232],
     pgate_l[233], pgate_l[234], pgate_l[235], pgate_l[236],
     pgate_l[237], pgate_l[238], pgate_l[239], pgate_l[240],
     pgate_l[241], pgate_l[242], pgate_l[243], pgate_l[244],
     pgate_l[245], pgate_l[246], pgate_l[247], pgate_l[248],
     pgate_l[249], pgate_l[250], pgate_l[251], pgate_l[252],
     pgate_l[253], pgate_l[254], pgate_l[255], pgate_l[256],
     pgate_l[257], pgate_l[258], pgate_l[259], pgate_l[260],
     pgate_l[261], pgate_l[262], pgate_l[263], pgate_l[264],
     pgate_l[265], pgate_l[266], pgate_l[267], pgate_l[268],
     pgate_l[269], pgate_l[270], pgate_l[271], pgate_l[272],
     pgate_l[273], pgate_l[274], pgate_l[275], pgate_l[276],
     pgate_l[277], pgate_l[278], pgate_l[279], pgate_l[280],
     pgate_l[281], pgate_l[282], pgate_l[283], pgate_l[284],
     pgate_l[285], pgate_l[286], pgate_l[287]}),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu1_b),
     .smc_write(smc_write_rowu1), .smc_rsr_inc(smc_row_inc_rowu1),
     .rsr_rst(smc_rsr_rst_rowu1), .por_rst(core_por_b_rowu1),
     .cram_wl_en(cram_wl_en_rowu1), .cram_vddoff(cram_vddoff_rowu1),
     .cram_rst(cram_rst_rowu1), .cram_pgateoff(cram_pgateoff_rowu1),
     .banksel(cm_banksel_bltld3_1_), .last_rsr(last_rsr[1]),
     .trst_b(trst_rowu1), .jtag_rowtest_rst(row_test_rowu1),
     .jtag_clk(tck_pad_rowu1));
ml_rowdrv_bank_1k Irowbl ( .vddctrl(vdd_cntl_l[143:0]),
     .wl(wl_l[143:0]), .reset(reset_l[143:0]), .pgate(pgate_l[143:0]),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu0_b),
     .smc_write(smc_write_rowu0), .smc_rsr_inc(smc_row_inc_rowu0),
     .rsr_rst(smc_rsr_rst_rowu0), .por_rst(core_por_b_rowu0),
     .cram_wl_en(cram_wl_en_rowu0), .cram_vddoff(cram_vddoff_rowu0),
     .cram_rst(cram_rst_rowu0), .cram_pgateoff(cram_pgateoff_rowu0),
     .banksel(cm_banksel_blbld1[0]), .last_rsr(last_rsr[0]),
     .trst_b(trst_rowu0), .jtag_rowtest_rst(row_test_rowu0),
     .jtag_clk(tck_pad_rowu0));
tielo I451_1_ ( .tielo(net129[0]));
tielo I451_0_ ( .tielo(net129[1]));
tielo I452 ( .tielo(net130));
sg_dffbuf_modified I261_1_ ( .r(net129[0]), .dffout(dff_out[1]),
     .d(cm_sdo_u1d[1]), .clk(net176));
sg_dffbuf_modified I261_0_ ( .r(net129[1]), .dffout(dff_out[0]),
     .d(cm_sdo_u1d[0]), .clk(net176));
sg_dffbuf_modified I289 ( .r(net130), .d(last_rsr[0]), .clk(net174),
     .dffout(last_rsr0));
bram_bufferx16 I381 ( .in(j_rst_bl1), .out(trst_rowu0));
bram_bufferx16 I391 ( .in(j_rst_bl2), .out(trst_rowu1));
bram_bufferx16 I392 ( .in(row_testl3), .out(row_test_rowu1));
bram_bufferx16 I393 ( .in(cram_pgateoffl2), .out(cram_pgateoff_rowu1));
bram_bufferx16 I394 ( .in(cram_rstl2), .out(cram_rst_rowu1));
bram_bufferx16 I395 ( .in(cram_wl_enl2), .out(cram_wl_en_rowu1));
bram_bufferx16 I396 ( .in(smc_writel2), .out(smc_write_rowu1));
bram_bufferx16 I397 ( .in(cram_vddoffl2), .out(cram_vddoff_rowu1));
bram_bufferx16 I398 ( .in(smc_row_incl2), .out(smc_row_inc_rowu1));
bram_bufferx16 I400 ( .in(smc_rsr_rstl2), .out(smc_rsr_rst_rowu1));
bram_bufferx16 I390 ( .in(smc_rsr_rstl1), .out(smc_rsr_rst_rowu0));
bram_bufferx16 I435 ( .in(tck_padl2), .out(tck_pad_rowu1));
bram_bufferx16 I384 ( .in(cram_rstl1), .out(cram_rst_rowu0));
bram_bufferx16 I290 ( .in(cm_clk_blbld), .out(net174));
bram_bufferx16 I260 ( .in(cm_clk_blbld), .out(net176));
bram_bufferx16 I385 ( .in(cram_vddoffl1), .out(cram_vddoff_rowu0));
bram_bufferx16 I386 ( .in(cram_wl_enl1), .out(cram_wl_en_rowu0));
bram_bufferx16 I387 ( .in(smc_row_incl1), .out(smc_row_inc_rowu0));
bram_bufferx16 I388 ( .in(smc_writel1), .out(smc_write_rowu0));
bram_bufferx16 I389 ( .in(core_por_bbl1), .out(core_por_b_rowu0));
bram_bufferx16 I383 ( .in(cram_pgateoffl1), .out(cram_pgateoff_rowu0));
bram_bufferx16 I437 ( .in(tck_padl1), .out(tck_pad_rowu0));
bram_bufferx16 I382 ( .in(row_testl2), .out(row_test_rowu0));
sg_bufx10 I421 ( .in(cf_lbank[479]), .out(monitor_celld[1]));
sg_bufx10 I235 ( .in(data_muxsel_bltld), .out(data_muxsel_bltld3));
sg_bufx10 I425 ( .in(monitor_celld[1]), .out(monitor_celld1[1]));
sg_bufx10 I424 ( .in(cf_lbank[300]), .out(monitor_celld2[0]));
sg_bufx10 I426 ( .in(monitor_celld1[1]), .out(monitor_celld2[1]));
sg_bufx10 I450_1_ ( .in(dff_out[1]), .out(cm_sdo_u1d1[1]));
sg_bufx10 I450_0_ ( .in(dff_out[0]), .out(cm_sdo_u1d1[0]));
sg_bufx10 I106_1_ ( .in(cm_sdo_u1[1]), .out(cm_sdo_u1d0[1]));
sg_bufx10 I106_0_ ( .in(cm_sdo_u1[0]), .out(cm_sdo_u1d0[0]));
sg_bufx10 I337 ( .in(core_por_bbl0), .out(core_por_bbl1));
sg_bufx10 I338 ( .in(smc_rsr_rstl0), .out(smc_rsr_rstl1));
sg_bufx10 I339 ( .in(row_testl1), .out(row_testl2));
sg_bufx10 I340 ( .in(j_rst_bl0), .out(j_rst_bl1));
sg_bufx10 I342 ( .in(smc_writel0), .out(smc_writel1));
sg_bufx10 I343 ( .in(smc_row_incl0), .out(smc_row_incl1));
sg_bufx10 I344 ( .in(cram_wl_enl0), .out(cram_wl_enl1));
sg_bufx10 I345 ( .in(cram_vddoffl0), .out(cram_vddoffl1));
sg_bufx10 I346 ( .in(cram_rstl0), .out(cram_rstl1));
sg_bufx10 I347 ( .in(cram_pgateoffl0), .out(cram_pgateoffl1));
sg_bufx10 I355 ( .in(cram_pgateoffl1), .out(cram_pgateoffl2));
sg_bufx10 I438 ( .in(tck_padl0), .out(tck_padl1));
sg_bufx10 I237 ( .in(data_muxsel1_bltld), .out(data_muxsel1_bltld3));
sg_bufx10 I351 ( .in(smc_row_incl1), .out(smc_row_incl2));
sg_bufx10 I368 ( .in(cram_pullup_bltld), .out(cram_pullup_bltld3));
sg_bufx10 I277 ( .in(cm_banksel_blbld[1]), .out(cm_banksel_bltld[1]));
sg_bufx10 I348 ( .in(smc_rsr_rstl1), .out(smc_rsr_rstl2));
sg_bufx10 I278_1_ ( .in(cm_sdo_u1d0[1]), .out(cm_sdo_u1d[1]));
sg_bufx10 I278_0_ ( .in(cm_sdo_u1d0[0]), .out(cm_sdo_u1d[0]));
sg_bufx10 I354 ( .in(cram_rstl1), .out(cram_rstl2));
sg_bufx10 I271 ( .in(data_muxsel1_blbld), .out(data_muxsel1_bltld));
sg_bufx10 I275 ( .in(cram_prec_blbld), .out(cram_prec_bltld));
sg_bufx10 I241 ( .in(en_8bconfig_b_bltld), .out(en_8bconfig_b_bltld3));
sg_bufx10 I353 ( .in(cram_vddoffl1), .out(cram_vddoffl2));
sg_bufx10 I357 ( .in(j_rst_bl1), .out(j_rst_bl2));
sg_bufx10 I356 ( .in(row_testl2), .out(row_testl3));
sg_bufx10 I273 ( .in(smc_wdis_dclk_blbld), .out(smc_wdis_dclk_bltld));
sg_bufx10 I279_1_ ( .in(cm_sdi_u1d[1]), .out(cm_sdi_u1d0[1]));
sg_bufx10 I279_0_ ( .in(cm_sdi_u1d[0]), .out(cm_sdi_u1d0[0]));
sg_bufx10 I272 ( .in(en_8bconfig_b_blbld), .out(en_8bconfig_b_bltld));
sg_bufx10 I274 ( .in(cram_write_blbld), .out(cram_write_bltld));
sg_bufx10 I239 ( .in(smc_wdis_dclk_bltld), .out(smc_wdis_dclk_bltld3));
sg_bufx10 I270 ( .in(data_muxsel_blbld), .out(data_muxsel_bltld));
sg_bufx10 I240 ( .in(cram_write_bltld), .out(cram_write_bltld3));
sg_bufx10 I238 ( .in(cram_prec_bltld), .out(cram_prec_bltld3));
sg_bufx10 I242 ( .in(cm_clk_bltld), .out(cm_clk_bltld3));
sg_bufx10 I236 ( .in(cm_banksel_bltld[1]), .out(cm_banksel_bltld3_1_));
sg_bufx10 I276 ( .in(cm_clk_blbld), .out(cm_clk_bltld));
sg_bufx10 I352 ( .in(cram_wl_enl1), .out(cram_wl_enl2));
sg_bufx10 I280_1_ ( .in(cm_sdi_u1d0[1]), .out(cm_sdi_u1d3[1]));
sg_bufx10 I280_0_ ( .in(cm_sdi_u1d0[0]), .out(cm_sdi_u1d3[0]));
sg_bufx10 I350 ( .in(smc_writel1), .out(smc_writel2));
sg_bufx10 I349 ( .in(core_por_bbl1), .out(core_por_b_rowu1));
sg_bufx10 I369 ( .in(cram_pullup_blbld), .out(cram_pullup_bltld));
sg_bufx10 I436 ( .in(tck_padl1), .out(tck_padl2));

endmodule
// Library - chip, Cell - CHIP_route_right1f, View - schematic
// LAST TIME SAVED: Jun 16 09:08:14 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module CHIP_route_right1f ( cm_banksel_bltld3_1_, cm_clk_bltld3,
     cm_sdi_u1d3[1:0], cm_sdo_u1d1[1:0], core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, last_rsr[1:0],
     monitor_celld2[1:0], pgate_r[287:0], reset_r[287:0],
     smc_wdis_dclk_bltld3, vdd_cntl_r[287:0], wl_r[287:0],
     cf_lbank[300], cf_lbank[479], cm_banksel_blbld1[0],
     cm_banksel_blbld[1], cm_clk_blbld, cm_sdi_u1d[1:0],
     cm_sdo_u1[1:0], core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0 );
output  cm_banksel_bltld3_1_, cm_clk_bltld3, core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, smc_wdis_dclk_bltld3;

input  cm_clk_blbld, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;

output [1:0]  cm_sdo_u1d1;
output [1:0]  cm_sdi_u1d3;
output [287:0]  pgate_r;
output [1:0]  last_rsr;
output [287:0]  vdd_cntl_r;
output [1:0]  monitor_celld2;
output [287:0]  reset_r;
output [287:0]  wl_r;

input [1:0]  cm_sdi_u1d;
input [0:0]  cm_banksel_blbld1;
input [300:479]  cf_lbank;
input [1:0]  cm_sdo_u1;
input [1:1]  cm_banksel_blbld;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u1d;

wire  [0:1]  net129;

wire  [1:0]  dff_out;

wire  [1:0]  cm_sdi_u1d0;

wire  [1:1]  cm_banksel_bltld;

wire  [1:1]  monitor_celld1;

wire  [1:0]  cm_sdo_u1d0;

wire  [1:1]  monitor_celld;



ml_rowdrv_bank_1k Irowul ( .vddctrl({vdd_cntl_r[144], vdd_cntl_r[145],
     vdd_cntl_r[146], vdd_cntl_r[147], vdd_cntl_r[148],
     vdd_cntl_r[149], vdd_cntl_r[150], vdd_cntl_r[151],
     vdd_cntl_r[152], vdd_cntl_r[153], vdd_cntl_r[154],
     vdd_cntl_r[155], vdd_cntl_r[156], vdd_cntl_r[157],
     vdd_cntl_r[158], vdd_cntl_r[159], vdd_cntl_r[160],
     vdd_cntl_r[161], vdd_cntl_r[162], vdd_cntl_r[163],
     vdd_cntl_r[164], vdd_cntl_r[165], vdd_cntl_r[166],
     vdd_cntl_r[167], vdd_cntl_r[168], vdd_cntl_r[169],
     vdd_cntl_r[170], vdd_cntl_r[171], vdd_cntl_r[172],
     vdd_cntl_r[173], vdd_cntl_r[174], vdd_cntl_r[175],
     vdd_cntl_r[176], vdd_cntl_r[177], vdd_cntl_r[178],
     vdd_cntl_r[179], vdd_cntl_r[180], vdd_cntl_r[181],
     vdd_cntl_r[182], vdd_cntl_r[183], vdd_cntl_r[184],
     vdd_cntl_r[185], vdd_cntl_r[186], vdd_cntl_r[187],
     vdd_cntl_r[188], vdd_cntl_r[189], vdd_cntl_r[190],
     vdd_cntl_r[191], vdd_cntl_r[192], vdd_cntl_r[193],
     vdd_cntl_r[194], vdd_cntl_r[195], vdd_cntl_r[196],
     vdd_cntl_r[197], vdd_cntl_r[198], vdd_cntl_r[199],
     vdd_cntl_r[200], vdd_cntl_r[201], vdd_cntl_r[202],
     vdd_cntl_r[203], vdd_cntl_r[204], vdd_cntl_r[205],
     vdd_cntl_r[206], vdd_cntl_r[207], vdd_cntl_r[208],
     vdd_cntl_r[209], vdd_cntl_r[210], vdd_cntl_r[211],
     vdd_cntl_r[212], vdd_cntl_r[213], vdd_cntl_r[214],
     vdd_cntl_r[215], vdd_cntl_r[216], vdd_cntl_r[217],
     vdd_cntl_r[218], vdd_cntl_r[219], vdd_cntl_r[220],
     vdd_cntl_r[221], vdd_cntl_r[222], vdd_cntl_r[223],
     vdd_cntl_r[224], vdd_cntl_r[225], vdd_cntl_r[226],
     vdd_cntl_r[227], vdd_cntl_r[228], vdd_cntl_r[229],
     vdd_cntl_r[230], vdd_cntl_r[231], vdd_cntl_r[232],
     vdd_cntl_r[233], vdd_cntl_r[234], vdd_cntl_r[235],
     vdd_cntl_r[236], vdd_cntl_r[237], vdd_cntl_r[238],
     vdd_cntl_r[239], vdd_cntl_r[240], vdd_cntl_r[241],
     vdd_cntl_r[242], vdd_cntl_r[243], vdd_cntl_r[244],
     vdd_cntl_r[245], vdd_cntl_r[246], vdd_cntl_r[247],
     vdd_cntl_r[248], vdd_cntl_r[249], vdd_cntl_r[250],
     vdd_cntl_r[251], vdd_cntl_r[252], vdd_cntl_r[253],
     vdd_cntl_r[254], vdd_cntl_r[255], vdd_cntl_r[256],
     vdd_cntl_r[257], vdd_cntl_r[258], vdd_cntl_r[259],
     vdd_cntl_r[260], vdd_cntl_r[261], vdd_cntl_r[262],
     vdd_cntl_r[263], vdd_cntl_r[264], vdd_cntl_r[265],
     vdd_cntl_r[266], vdd_cntl_r[267], vdd_cntl_r[268],
     vdd_cntl_r[269], vdd_cntl_r[270], vdd_cntl_r[271],
     vdd_cntl_r[272], vdd_cntl_r[273], vdd_cntl_r[274],
     vdd_cntl_r[275], vdd_cntl_r[276], vdd_cntl_r[277],
     vdd_cntl_r[278], vdd_cntl_r[279], vdd_cntl_r[280],
     vdd_cntl_r[281], vdd_cntl_r[282], vdd_cntl_r[283],
     vdd_cntl_r[284], vdd_cntl_r[285], vdd_cntl_r[286],
     vdd_cntl_r[287]}), .wl({wl_r[144], wl_r[145], wl_r[146],
     wl_r[147], wl_r[148], wl_r[149], wl_r[150], wl_r[151], wl_r[152],
     wl_r[153], wl_r[154], wl_r[155], wl_r[156], wl_r[157], wl_r[158],
     wl_r[159], wl_r[160], wl_r[161], wl_r[162], wl_r[163], wl_r[164],
     wl_r[165], wl_r[166], wl_r[167], wl_r[168], wl_r[169], wl_r[170],
     wl_r[171], wl_r[172], wl_r[173], wl_r[174], wl_r[175], wl_r[176],
     wl_r[177], wl_r[178], wl_r[179], wl_r[180], wl_r[181], wl_r[182],
     wl_r[183], wl_r[184], wl_r[185], wl_r[186], wl_r[187], wl_r[188],
     wl_r[189], wl_r[190], wl_r[191], wl_r[192], wl_r[193], wl_r[194],
     wl_r[195], wl_r[196], wl_r[197], wl_r[198], wl_r[199], wl_r[200],
     wl_r[201], wl_r[202], wl_r[203], wl_r[204], wl_r[205], wl_r[206],
     wl_r[207], wl_r[208], wl_r[209], wl_r[210], wl_r[211], wl_r[212],
     wl_r[213], wl_r[214], wl_r[215], wl_r[216], wl_r[217], wl_r[218],
     wl_r[219], wl_r[220], wl_r[221], wl_r[222], wl_r[223], wl_r[224],
     wl_r[225], wl_r[226], wl_r[227], wl_r[228], wl_r[229], wl_r[230],
     wl_r[231], wl_r[232], wl_r[233], wl_r[234], wl_r[235], wl_r[236],
     wl_r[237], wl_r[238], wl_r[239], wl_r[240], wl_r[241], wl_r[242],
     wl_r[243], wl_r[244], wl_r[245], wl_r[246], wl_r[247], wl_r[248],
     wl_r[249], wl_r[250], wl_r[251], wl_r[252], wl_r[253], wl_r[254],
     wl_r[255], wl_r[256], wl_r[257], wl_r[258], wl_r[259], wl_r[260],
     wl_r[261], wl_r[262], wl_r[263], wl_r[264], wl_r[265], wl_r[266],
     wl_r[267], wl_r[268], wl_r[269], wl_r[270], wl_r[271], wl_r[272],
     wl_r[273], wl_r[274], wl_r[275], wl_r[276], wl_r[277], wl_r[278],
     wl_r[279], wl_r[280], wl_r[281], wl_r[282], wl_r[283], wl_r[284],
     wl_r[285], wl_r[286], wl_r[287]}), .reset({reset_r[144],
     reset_r[145], reset_r[146], reset_r[147], reset_r[148],
     reset_r[149], reset_r[150], reset_r[151], reset_r[152],
     reset_r[153], reset_r[154], reset_r[155], reset_r[156],
     reset_r[157], reset_r[158], reset_r[159], reset_r[160],
     reset_r[161], reset_r[162], reset_r[163], reset_r[164],
     reset_r[165], reset_r[166], reset_r[167], reset_r[168],
     reset_r[169], reset_r[170], reset_r[171], reset_r[172],
     reset_r[173], reset_r[174], reset_r[175], reset_r[176],
     reset_r[177], reset_r[178], reset_r[179], reset_r[180],
     reset_r[181], reset_r[182], reset_r[183], reset_r[184],
     reset_r[185], reset_r[186], reset_r[187], reset_r[188],
     reset_r[189], reset_r[190], reset_r[191], reset_r[192],
     reset_r[193], reset_r[194], reset_r[195], reset_r[196],
     reset_r[197], reset_r[198], reset_r[199], reset_r[200],
     reset_r[201], reset_r[202], reset_r[203], reset_r[204],
     reset_r[205], reset_r[206], reset_r[207], reset_r[208],
     reset_r[209], reset_r[210], reset_r[211], reset_r[212],
     reset_r[213], reset_r[214], reset_r[215], reset_r[216],
     reset_r[217], reset_r[218], reset_r[219], reset_r[220],
     reset_r[221], reset_r[222], reset_r[223], reset_r[224],
     reset_r[225], reset_r[226], reset_r[227], reset_r[228],
     reset_r[229], reset_r[230], reset_r[231], reset_r[232],
     reset_r[233], reset_r[234], reset_r[235], reset_r[236],
     reset_r[237], reset_r[238], reset_r[239], reset_r[240],
     reset_r[241], reset_r[242], reset_r[243], reset_r[244],
     reset_r[245], reset_r[246], reset_r[247], reset_r[248],
     reset_r[249], reset_r[250], reset_r[251], reset_r[252],
     reset_r[253], reset_r[254], reset_r[255], reset_r[256],
     reset_r[257], reset_r[258], reset_r[259], reset_r[260],
     reset_r[261], reset_r[262], reset_r[263], reset_r[264],
     reset_r[265], reset_r[266], reset_r[267], reset_r[268],
     reset_r[269], reset_r[270], reset_r[271], reset_r[272],
     reset_r[273], reset_r[274], reset_r[275], reset_r[276],
     reset_r[277], reset_r[278], reset_r[279], reset_r[280],
     reset_r[281], reset_r[282], reset_r[283], reset_r[284],
     reset_r[285], reset_r[286], reset_r[287]}), .pgate({pgate_r[144],
     pgate_r[145], pgate_r[146], pgate_r[147], pgate_r[148],
     pgate_r[149], pgate_r[150], pgate_r[151], pgate_r[152],
     pgate_r[153], pgate_r[154], pgate_r[155], pgate_r[156],
     pgate_r[157], pgate_r[158], pgate_r[159], pgate_r[160],
     pgate_r[161], pgate_r[162], pgate_r[163], pgate_r[164],
     pgate_r[165], pgate_r[166], pgate_r[167], pgate_r[168],
     pgate_r[169], pgate_r[170], pgate_r[171], pgate_r[172],
     pgate_r[173], pgate_r[174], pgate_r[175], pgate_r[176],
     pgate_r[177], pgate_r[178], pgate_r[179], pgate_r[180],
     pgate_r[181], pgate_r[182], pgate_r[183], pgate_r[184],
     pgate_r[185], pgate_r[186], pgate_r[187], pgate_r[188],
     pgate_r[189], pgate_r[190], pgate_r[191], pgate_r[192],
     pgate_r[193], pgate_r[194], pgate_r[195], pgate_r[196],
     pgate_r[197], pgate_r[198], pgate_r[199], pgate_r[200],
     pgate_r[201], pgate_r[202], pgate_r[203], pgate_r[204],
     pgate_r[205], pgate_r[206], pgate_r[207], pgate_r[208],
     pgate_r[209], pgate_r[210], pgate_r[211], pgate_r[212],
     pgate_r[213], pgate_r[214], pgate_r[215], pgate_r[216],
     pgate_r[217], pgate_r[218], pgate_r[219], pgate_r[220],
     pgate_r[221], pgate_r[222], pgate_r[223], pgate_r[224],
     pgate_r[225], pgate_r[226], pgate_r[227], pgate_r[228],
     pgate_r[229], pgate_r[230], pgate_r[231], pgate_r[232],
     pgate_r[233], pgate_r[234], pgate_r[235], pgate_r[236],
     pgate_r[237], pgate_r[238], pgate_r[239], pgate_r[240],
     pgate_r[241], pgate_r[242], pgate_r[243], pgate_r[244],
     pgate_r[245], pgate_r[246], pgate_r[247], pgate_r[248],
     pgate_r[249], pgate_r[250], pgate_r[251], pgate_r[252],
     pgate_r[253], pgate_r[254], pgate_r[255], pgate_r[256],
     pgate_r[257], pgate_r[258], pgate_r[259], pgate_r[260],
     pgate_r[261], pgate_r[262], pgate_r[263], pgate_r[264],
     pgate_r[265], pgate_r[266], pgate_r[267], pgate_r[268],
     pgate_r[269], pgate_r[270], pgate_r[271], pgate_r[272],
     pgate_r[273], pgate_r[274], pgate_r[275], pgate_r[276],
     pgate_r[277], pgate_r[278], pgate_r[279], pgate_r[280],
     pgate_r[281], pgate_r[282], pgate_r[283], pgate_r[284],
     pgate_r[285], pgate_r[286], pgate_r[287]}),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu1_b),
     .smc_write(smc_write_rowu1), .smc_rsr_inc(smc_row_inc_rowu1),
     .rsr_rst(smc_rsr_rst_rowu1), .por_rst(core_por_b_rowu1),
     .cram_wl_en(cram_wl_en_rowu1), .cram_vddoff(cram_vddoff_rowu1),
     .cram_rst(cram_rst_rowu1), .cram_pgateoff(cram_pgateoff_rowu1),
     .banksel(cm_banksel_bltld3_1_), .last_rsr(last_rsr[1]),
     .trst_b(trst_rowu1), .jtag_rowtest_rst(row_test_rowu1),
     .jtag_clk(tck_pad_rowu1));
ml_rowdrv_bank_1k Irowbl ( .vddctrl(vdd_cntl_r[143:0]),
     .wl(wl_r[143:0]), .reset(reset_r[143:0]), .pgate(pgate_r[143:0]),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu0_b),
     .smc_write(smc_write_rowu0), .smc_rsr_inc(smc_row_inc_rowu0),
     .rsr_rst(smc_rsr_rst_rowu0), .por_rst(core_por_b_rowu0),
     .cram_wl_en(cram_wl_en_rowu0), .cram_vddoff(cram_vddoff_rowu0),
     .cram_rst(cram_rst_rowu0), .cram_pgateoff(cram_pgateoff_rowu0),
     .banksel(cm_banksel_blbld1[0]), .last_rsr(last_rsr[0]),
     .trst_b(trst_rowu0), .jtag_rowtest_rst(row_test_rowu0),
     .jtag_clk(tck_pad_rowu0));
tielo I5_1_ ( .tielo(net129[0]));
tielo I5_0_ ( .tielo(net129[1]));
tielo I4 ( .tielo(net130));
sg_dffbuf_modified I70_1_ ( .r(net129[0]), .dffout(dff_out[1]),
     .d(cm_sdo_u1d[1]), .clk(net176));
sg_dffbuf_modified I70_0_ ( .r(net129[1]), .dffout(dff_out[0]),
     .d(cm_sdo_u1d[0]), .clk(net176));
sg_dffbuf_modified I57 ( .r(net130), .d(last_rsr[0]), .clk(net174),
     .dffout(last_rsr0));
bram_bufferx16 I33 ( .in(j_rst_bl1), .out(trst_rowu0));
bram_bufferx16 I23 ( .in(j_rst_bl2), .out(trst_rowu1));
bram_bufferx16 I22 ( .in(row_testl3), .out(row_test_rowu1));
bram_bufferx16 I21 ( .in(cram_pgateoffl2), .out(cram_pgateoff_rowu1));
bram_bufferx16 I20 ( .in(cram_rstl2), .out(cram_rst_rowu1));
bram_bufferx16 I19 ( .in(cram_wl_enl2), .out(cram_wl_en_rowu1));
bram_bufferx16 I18 ( .in(smc_writel2), .out(smc_write_rowu1));
bram_bufferx16 I17 ( .in(cram_vddoffl2), .out(cram_vddoff_rowu1));
bram_bufferx16 I16 ( .in(smc_row_incl2), .out(smc_row_inc_rowu1));
bram_bufferx16 I15 ( .in(smc_rsr_rstl2), .out(smc_rsr_rst_rowu1));
bram_bufferx16 I24 ( .in(smc_rsr_rstl1), .out(smc_rsr_rst_rowu0));
bram_bufferx16 I10 ( .in(tck_padl2), .out(tck_pad_rowu1));
bram_bufferx16 I30 ( .in(cram_rstl1), .out(cram_rst_rowu0));
bram_bufferx16 I56 ( .in(cm_clk_blbld), .out(net174));
bram_bufferx16 I71 ( .in(cm_clk_blbld), .out(net176));
bram_bufferx16 I29 ( .in(cram_vddoffl1), .out(cram_vddoff_rowu0));
bram_bufferx16 I28 ( .in(cram_wl_enl1), .out(cram_wl_en_rowu0));
bram_bufferx16 I27 ( .in(smc_row_incl1), .out(smc_row_inc_rowu0));
bram_bufferx16 I26 ( .in(smc_writel1), .out(smc_write_rowu0));
bram_bufferx16 I25 ( .in(core_por_bbl1), .out(core_por_b_rowu0));
bram_bufferx16 I31 ( .in(cram_pgateoffl1), .out(cram_pgateoff_rowu0));
bram_bufferx16 I8 ( .in(tck_padl1), .out(tck_pad_rowu0));
bram_bufferx16 I32 ( .in(row_testl2), .out(row_test_rowu0));
sg_bufx10 I14 ( .in(cf_lbank[479]), .out(monitor_celld[1]));
sg_bufx10 I79 ( .in(data_muxsel_bltld), .out(data_muxsel_bltld3));
sg_bufx10 I12 ( .in(monitor_celld[1]), .out(monitor_celld1[1]));
sg_bufx10 I13 ( .in(cf_lbank[300]), .out(monitor_celld2[0]));
sg_bufx10 I11 ( .in(monitor_celld1[1]), .out(monitor_celld2[1]));
sg_bufx10 I6_1_ ( .in(dff_out[1]), .out(cm_sdo_u1d1[1]));
sg_bufx10 I6_0_ ( .in(dff_out[0]), .out(cm_sdo_u1d1[0]));
sg_bufx10 I80_1_ ( .in(cm_sdo_u1[1]), .out(cm_sdo_u1d0[1]));
sg_bufx10 I80_0_ ( .in(cm_sdo_u1[0]), .out(cm_sdo_u1d0[0]));
sg_bufx10 I55 ( .in(core_por_bbl0), .out(core_por_bbl1));
sg_bufx10 I54 ( .in(smc_rsr_rstl0), .out(smc_rsr_rstl1));
sg_bufx10 I53 ( .in(row_testl1), .out(row_testl2));
sg_bufx10 I52 ( .in(j_rst_bl0), .out(j_rst_bl1));
sg_bufx10 I51 ( .in(smc_writel0), .out(smc_writel1));
sg_bufx10 I50 ( .in(smc_row_incl0), .out(smc_row_incl1));
sg_bufx10 I49 ( .in(cram_wl_enl0), .out(cram_wl_enl1));
sg_bufx10 I48 ( .in(cram_vddoffl0), .out(cram_vddoffl1));
sg_bufx10 I47 ( .in(cram_rstl0), .out(cram_rstl1));
sg_bufx10 I46 ( .in(cram_pgateoffl0), .out(cram_pgateoffl1));
sg_bufx10 I38 ( .in(cram_pgateoffl1), .out(cram_pgateoffl2));
sg_bufx10 I7 ( .in(tck_padl0), .out(tck_padl1));
sg_bufx10 I77 ( .in(data_muxsel1_bltld), .out(data_muxsel1_bltld3));
sg_bufx10 I42 ( .in(smc_row_incl1), .out(smc_row_incl2));
sg_bufx10 I35 ( .in(cram_pullup_bltld), .out(cram_pullup_bltld3));
sg_bufx10 I61 ( .in(cm_banksel_blbld[1]), .out(cm_banksel_bltld[1]));
sg_bufx10 I45 ( .in(smc_rsr_rstl1), .out(smc_rsr_rstl2));
sg_bufx10 I60_1_ ( .in(cm_sdo_u1d0[1]), .out(cm_sdo_u1d[1]));
sg_bufx10 I60_0_ ( .in(cm_sdo_u1d0[0]), .out(cm_sdo_u1d[0]));
sg_bufx10 I39 ( .in(cram_rstl1), .out(cram_rstl2));
sg_bufx10 I68 ( .in(data_muxsel1_blbld), .out(data_muxsel1_bltld));
sg_bufx10 I63 ( .in(cram_prec_blbld), .out(cram_prec_bltld));
sg_bufx10 I73 ( .in(en_8bconfig_b_bltld), .out(en_8bconfig_b_bltld3));
sg_bufx10 I40 ( .in(cram_vddoffl1), .out(cram_vddoffl2));
sg_bufx10 I36 ( .in(j_rst_bl1), .out(j_rst_bl2));
sg_bufx10 I37 ( .in(row_testl2), .out(row_testl3));
sg_bufx10 I65 ( .in(smc_wdis_dclk_blbld), .out(smc_wdis_dclk_bltld));
sg_bufx10 I59_1_ ( .in(cm_sdi_u1d[1]), .out(cm_sdi_u1d0[1]));
sg_bufx10 I59_0_ ( .in(cm_sdi_u1d[0]), .out(cm_sdi_u1d0[0]));
sg_bufx10 I67 ( .in(en_8bconfig_b_blbld), .out(en_8bconfig_b_bltld));
sg_bufx10 I64 ( .in(cram_write_blbld), .out(cram_write_bltld));
sg_bufx10 I75 ( .in(smc_wdis_dclk_bltld), .out(smc_wdis_dclk_bltld3));
sg_bufx10 I69 ( .in(data_muxsel_blbld), .out(data_muxsel_bltld));
sg_bufx10 I74 ( .in(cram_write_bltld), .out(cram_write_bltld3));
sg_bufx10 I76 ( .in(cram_prec_bltld), .out(cram_prec_bltld3));
sg_bufx10 I72 ( .in(cm_clk_bltld), .out(cm_clk_bltld3));
sg_bufx10 I78 ( .in(cm_banksel_bltld[1]), .out(cm_banksel_bltld3_1_));
sg_bufx10 I62 ( .in(cm_clk_blbld), .out(cm_clk_bltld));
sg_bufx10 I41 ( .in(cram_wl_enl1), .out(cram_wl_enl2));
sg_bufx10 I58_1_ ( .in(cm_sdi_u1d0[1]), .out(cm_sdi_u1d3[1]));
sg_bufx10 I58_0_ ( .in(cm_sdi_u1d0[0]), .out(cm_sdi_u1d3[0]));
sg_bufx10 I43 ( .in(smc_writel1), .out(smc_writel2));
sg_bufx10 I44 ( .in(core_por_bbl1), .out(core_por_b_rowu1));
sg_bufx10 I34 ( .in(cram_pullup_blbld), .out(cram_pullup_bltld));
sg_bufx10 I9 ( .in(tck_padl1), .out(tck_padl2));

endmodule
// Library - leafcell, Cell - fabric_buf8k, View - schematic
// LAST TIME SAVED: Jan 15 15:42:13 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module fabric_buf8k ( f_out, f_in );
output  f_out;

input  f_in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I252 ( .A(net6), .Y(f_out));
inv_hvt I248 ( .A(f_in), .Y(net6));

endmodule
// Library - xpmem, Cell - ml_blsa_clk_buf, View - schematic
// LAST TIME SAVED: Sep  5 15:09:27 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_clk_buf ( o, in );
output  o;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_powersurg_buf, View - schematic
// LAST TIME SAVED: Jul 31 18:29:48 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_powersurg_buf ( o, in );
output  o;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I404 ( .A(net016), .Y(net012));
inv_hvt I405 ( .A(net012), .Y(o));
inv_hvt I391 ( .A(net77), .Y(net016));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_dff_bl, View - schematic
// LAST TIME SAVED: Jan 30 16:47:38 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_dff_bl ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - xpmem, Cell - ml_blsa_sch, View - schematic
// LAST TIME SAVED: Jan 30 16:47:19 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_sch ( dataout, bl, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, datain, latch_clock, latch_reset, smc_wdic_clk );
output  dataout;

inout  bl;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, datain,
     latch_clock, latch_reset, smc_wdic_clk;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff_bl Idff ( .R(latch_reset), .D(dff_in), .CLK(latch_clock),
     .QN(write_data_b), .Q(dff_data));
nor2_hvt I223 ( .A(net084), .B(write_data_b), .Y(n_gate));
inv_hvt I163 ( .A(write_data_b), .Y(dataout));
inv_hvt I159 ( .A(cram_prec), .Y(net0161));
inv_hvt I160 ( .A(cram_write), .Y(net084));
mux2_hvt I161 ( .in1(sa_out), .in0(datain), .out(latch_in),
     .sel(data_muxsel));
mux2_hvt I164 ( .in1(dff_data), .in0(latch_in), .out(dff_in),
     .sel(smc_wdic_clk));
nch_hvt  MN12 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN8 ( .D(sa_out), .B(gnd_), .G(cram_pullup_b), .S(gnd_));
nch_hvt  MN10 ( .D(net0166), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN13 ( .D(net0184), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN3 ( .D(sa_out), .B(gnd_), .G(bl), .S(gnd_));
nch_hvt  MN6 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
pch_hvt  MP8 ( .D(net0148), .B(vdd_), .G(dataout), .S(vdd_));
pch_hvt  MP9 ( .D(bl), .B(vdd_), .G(net084), .S(net0148));
pch_hvt  MP13 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP12 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP14 ( .D(net0208), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP4 ( .D(net0143), .B(vdd_), .G(cram_pullup_b), .S(vdd_));
pch_hvt  MP5 ( .D(sa_out), .B(vdd_), .G(bl), .S(net0143));
pch_hvt  MP15 ( .D(net0204), .B(vdd_), .G(net0161), .S(vdd_));

endmodule
// Library - xpmem, Cell - ml_blsa_tile, View - schematic
// LAST TIME SAVED: Sep  5 14:53:52 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_tile ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [53:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [53:0]  dataout;

wire  [13:0]  ck;



ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
inv_hvt I172 ( .A(net48), .Y(data_out));
inv_hvt I171 ( .A(dataout[53]), .Y(net48));
ml_powersurg_buf I161 ( .in(cram_write), .o(net53));
ml_powersurg_buf I165 ( .in(net57), .o(net55));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net57));
ml_powersurg_buf I163 ( .in(net55), .o(net59));
ml_powersurg_buf I162 ( .in(net65), .o(net61));
ml_powersurg_buf I169 ( .in(net61), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net53), .o(net65));
ml_powersurg_buf I168 ( .in(net59), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_47_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[47]),
     .dataout(dataout[47]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_46_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[46]),
     .dataout(dataout[46]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_45_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[45]),
     .dataout(dataout[45]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_44_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[44]),
     .dataout(dataout[44]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_43_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[43]),
     .dataout(dataout[43]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_42_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[42]),
     .dataout(dataout[42]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_41_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_40_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_39_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_38_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_37_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_36_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_35_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_34_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_33_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_32_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net55));
ml_blsa_sch I170_53_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[52]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[53]),
     .dataout(dataout[53]), .cram_prec(net57));
ml_blsa_sch I170_52_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[51]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[52]),
     .dataout(dataout[52]), .cram_prec(net57));
ml_blsa_sch I170_51_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[50]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[51]),
     .dataout(dataout[51]), .cram_prec(net57));
ml_blsa_sch I170_50_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[49]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[50]),
     .dataout(dataout[50]), .cram_prec(net57));
ml_blsa_sch I170_49_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[48]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[49]),
     .dataout(dataout[49]), .cram_prec(net57));
ml_blsa_sch I170_48_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[47]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[48]),
     .dataout(dataout[48]), .cram_prec(net57));
ml_blsa_sch Iml_blsa_sch_31_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_30_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_29_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_28_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_27_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_26_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_25_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_24_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_23_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_22_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_21_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_20_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_19_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_18_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net59));

endmodule
// Library - xpmem, Cell - ml_buf_ice5, View - schematic
// LAST TIME SAVED: Aug 13 13:53:01 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_buf_ice5 ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));
inv_hvt I391 ( .A(net77), .Y(o));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_last, View - schematic
// LAST TIME SAVED: Aug 28 08:58:43 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_tile_last ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [17:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [17:0]  dataout;

wire  [4:0]  ck;



tiehi I186 ( .tiehi(net040));
ml_dff_bl Idff ( .R(latch_reset), .D(dataout[16]), .CLK(ck[0]),
     .QN(net50), .Q(net45));
ml_dff_bl I179 ( .R(latch_reset), .D(net58), .CLK(ck[0]), .QN(net49),
     .Q(net61));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_buf_ice5 I205 ( .in(net61), .o(data_out), .sel(net040));
mux2_hvt I174 ( .in1(net45), .in0(dataout[17]), .out(net58),
     .sel(data_muxsel));
ml_powersurg_buf I169 ( .in(cram_write), .o(cram_write_out));
ml_powersurg_buf I168 ( .in(cram_prec), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[16]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[17]), .dataout(dataout[17]));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[15]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[16]), .dataout(dataout[16]));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));

endmodule
// Library - xpmem, Cell - ml_blprecwrt_en, View - schematic
// LAST TIME SAVED: May 16 10:09:58 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blprecwrt_en ( data_out, action, clkin, data_in, rst );
output  data_out;

input  action, clkin, data_in, rst;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I161 ( .A(net89), .Y(net88));
inv_hvt I162 ( .A(action), .Y(net86));
inv_hvt I165 ( .A(net98), .Y(data_out));
nand3_hvt I160 ( .Y(net89), .B(data_in), .C(action), .A(clkin));
nor2_hvt I385 ( .A(net88), .B(net94), .Y(net98));
nor3_hvt I387 ( .B(net86), .Y(net94), .A(net98), .C(rst));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex1_last, View - schematic
// LAST TIME SAVED: Jan 26 15:30:32 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_tilex1_last ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [71:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_0 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_dic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(datain_io), .cram_write_out(wrt_en_last),
     .cram_prec_out(prec_en_last), .bl(bl[53:0]));
ml_blsa_tile_last Iml_blsa_tile_last ( .bl(bl[71:54]),
     .latch_reset(latch_reset_buf), .datain(datain_io),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .latch_clock(latch_clock_out), .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_dic_clk_buf));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
inv_hvt I185 ( .A(smc_wdic_clk), .Y(net091));
inv_hvt I184 ( .A(net091), .Y(smc_dic_clk_buf));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex1, View - schematic
// LAST TIME SAVED: Jan 26 13:57:24 2009
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_tilex1 ( data_out, latch_clock_out, prec_out, wrt_out,
     bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [53:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_0 ( .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_last), .cram_prec_out(prec_en_last),
     .bl(bl[53:0]));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
inv_hvt I183 ( .A(net088), .Y(smc_wdic_clk_buf));
inv_hvt I184 ( .A(smc_wdic_clk), .Y(net088));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - misc, Cell - smc_and_jtag_ice8f, View - schematic
// LAST TIME SAVED: Aug  8 16:20:55 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module smc_and_jtag_ice8f ( bm_bank_sdi, bm_banksel, bm_clk, bm_init,
     bm_rcapmux_en, bm_sa, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_banksel, cm_clk, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2, cm_sdi_u3, data_muxsel, data_muxsel1,
     en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0, j_hiz_b,
     j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck, j_tdi,
     j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, psdo, rst_b,
     smc_load_nvcm_bstream, smc_osc_fsel, smc_oscoff_b, smc_podt_off,
     smc_podt_rst, smc_read, smc_row_inc, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rsr_rst, smc_rwl_en, smc_seq_rst,
     smc_wcram_rst, smc_wdis_dclk, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out_b, tdo_oe_pad, tdo_pad,
     bm_bank_sdo, boot, bp0, bschain_sdo, cdone_in, cm_last_rsr,
     cm_monitor_cell, cm_sdo_u0, cm_sdo_u1, cm_sdo_u2, cm_sdo_u3,
     cnt_podt_out, coldboot_sel, creset_b, idcode_msb20bits, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     osc_clk, por_b, psdi, spi_clk_in, spi_sdi, spi_ss_in_b, tck_pad,
     tdi_pad, tms_pad, trst_pad, warmboot_sel );
output  bm_clk, bm_init, bm_rcapmux_en, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_clk, data_muxsel,
     data_muxsel1, en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0,
     j_hiz_b, j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck,
     j_tdi, j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, rst_b,
     smc_load_nvcm_bstream, smc_oscoff_b, smc_podt_off, smc_podt_rst,
     smc_read, smc_row_inc, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rsr_rst, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_wdis_dclk, smc_write, smc_wset_prec, smc_wset_precgnd,
     smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_oe_pad, tdo_pad;

input  boot, bp0, bschain_sdo, cdone_in, cm_last_rsr, cnt_podt_out,
     creset_b, nvcm_boot, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, osc_clk, por_b, spi_clk_in, spi_sdi,
     spi_ss_in_b, tck_pad, tdi_pad, tms_pad, trst_pad;

output [3:0]  bm_bank_sdi;
output [3:0]  bm_banksel;
output [3:0]  cm_banksel;
output [1:0]  cm_sdi_u2;
output [1:0]  cm_sdi_u1;
output [7:1]  psdo;
output [1:0]  smc_osc_fsel;
output [7:0]  bm_sa;
output [1:0]  cm_sdi_u0;
output [1:0]  cm_sdi_u3;

input [3:0]  cm_monitor_cell;
input [1:0]  cm_sdo_u3;
input [1:0]  cm_sdo_u0;
input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdo_u2;
input [1:0]  warmboot_sel;
input [19:0]  idcode_msb20bits;
input [3:0]  bm_bank_sdo;
input [7:1]  psdi;
input [1:0]  coldboot_sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - xpmem, Cell - ml_blsa_tile_bram10k, View - schematic
// LAST TIME SAVED: Mar 20 10:20:41 2008
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_tile_bram10k ( cram_prec_out, cram_write_out, data_out,
     para_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, para_en, para_in,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out, para_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, para_en, para_in, smc_wdic_clk;

inout [41:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:4]  data_dummy_in;

wire  [0:41]  dataout;

wire  [0:14]  ck;

wire  [0:5]  data_in;



ml_dff_bl I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net97), .Q(net119));
ml_dff_bl I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net92), .Q(data_dummy_in[4]));
ml_dff_bl I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net87), .Q(data_dummy_in[2]));
ml_dff_bl I179 ( .R(latch_reset), .D(data_in[0]), .CLK(ck[14]),
     .QN(net82), .Q(data_dummy_in[1]));
ml_dff_bl I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net77), .Q(data_dummy_in[3]));
ml_blsa_clk_buf I192_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I192_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I192_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I192_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I192_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I192_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I192_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I192_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I192_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I192_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I192_0_ ( .in(latch_clock), .o(ck[0]));
mux2_hvt I194 ( .in1(data_dummy_in[2]), .in0(dataout[3]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I161 ( .in1(para_in), .in0(dataout[1]), .out(data_out_mux),
     .sel(para_en));
mux2_hvt I199 ( .in1(net119), .in0(dataout[6]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I198 ( .in1(data_dummy_in[4]), .in0(dataout[5]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I196 ( .in1(data_dummy_in[1]), .in0(dataout[2]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I197 ( .in1(data_dummy_in[3]), .in0(dataout[4]),
     .out(data_in[3]), .sel(data_muxsel1));
inv_hvt I262 ( .A(data_out_mux), .Y(net151));
inv_hvt I261 ( .A(net151), .Y(data_in[0]));
inv_hvt I175 ( .A(dataout[1]), .Y(net154));
inv_hvt I176 ( .A(net154), .Y(para_out));
inv_hvt I172 ( .A(net160), .Y(data_out));
inv_hvt I171 ( .A(dataout[41]), .Y(net160));
inv_hvt I200 ( .A(net133), .Y(net0132));
inv_hvt I201 ( .A(net0132), .Y(net0133));
inv_hvt I202 ( .A(net0133), .Y(net0131));
inv_hvt I229 ( .A(latch_clock), .Y(net133));
inv_hvt I203 ( .A(net0131), .Y(net0126));
inv_hvt I204 ( .A(net0126), .Y(ck[14]));
ml_powersurg_buf I165 ( .in(cram_prec), .o(net162));
ml_powersurg_buf I163 ( .in(net162), .o(net164));
ml_powersurg_buf I162 ( .in(net170), .o(net166));
ml_powersurg_buf I169 ( .in(net166), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(cram_write), .o(net170));
ml_powersurg_buf I168 ( .in(net164), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(data_in[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(data_in[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_41_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_40_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_39_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_38_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_37_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_36_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_35_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_34_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_33_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_32_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_31_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_30_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_29_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_28_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_27_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_26_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_25_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_24_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_23_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_22_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_21_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_20_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_19_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_18_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[14]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[15]),
     .dataout(dataout[15]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[13]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[14]),
     .dataout(dataout[14]), .cram_prec(net164));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_bram10k, View - schematic
// LAST TIME SAVED: Nov 30 09:32:34 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_tilex2_bram10k ( data_out, latch_clock_out, para_out,
     prec_out, wrt_out, bl, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, datain, latch_clock_in, latch_reset,
     para_en, para_in, prec_in, smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, para_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, para_en, para_in, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in;

inout [95:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile_bram10k Iml_blsa_tile_0 ( .para_en(para_en),
     .para_in(para_in), .para_out(para_out), .bl(bl[41:0]),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_en_last),
     .cram_prec_out(prec_en_last));
ml_blsa_tile Iml_blsa_tile_1 ( .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[95:42]));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
inv_hvt I183 ( .A(net088), .Y(smc_wdic_clk_buf));
inv_hvt I184 ( .A(smc_wdic_clk), .Y(net088));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_1st, View - schematic
// LAST TIME SAVED: Sep  6 14:29:58 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_tile_1st ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [55:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:4]  data_dummy_in;

wire  [1:5]  data_in;

wire  [0:55]  dataout;

wire  [0:14]  ck;



ml_dff_bl I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net132), .Q(net154));
ml_dff_bl I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net137), .Q(data_dummy_in[4]));
ml_dff_bl I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net142), .Q(data_dummy_in[2]));
ml_dff_bl I179 ( .R(latch_reset), .D(datain), .CLK(ck[14]),
     .QN(net147), .Q(data_dummy_in[1]));
ml_dff_bl I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net152), .Q(data_dummy_in[3]));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_blsa_sch Iml_blsa_sch_15_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[14]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_14_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[13]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_13_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[12]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_12_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[11]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_11_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[10]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_10_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[9]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_9_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[8]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_8_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[7]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_7_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[6]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_6_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_5_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_4_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[4]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_3_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[3]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_2_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[2]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_1_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[1]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_0_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(datain), .cram_prec(cram_prec_out),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_47_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[47]),
     .dataout(dataout[47]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_46_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[46]),
     .dataout(dataout[46]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_45_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[45]),
     .dataout(dataout[45]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_44_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[44]),
     .dataout(dataout[44]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_43_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[43]),
     .dataout(dataout[43]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_42_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[42]),
     .dataout(dataout[42]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_41_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[41]),
     .dataout(dataout[41]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_40_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[40]),
     .dataout(dataout[40]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_39_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[39]),
     .dataout(dataout[39]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_38_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[38]),
     .dataout(dataout[38]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_37_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[37]),
     .dataout(dataout[37]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_36_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[36]),
     .dataout(dataout[36]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_35_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[35]),
     .dataout(dataout[35]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_34_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[34]),
     .dataout(dataout[34]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_33_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[33]),
     .dataout(dataout[33]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_32_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[32]),
     .dataout(dataout[32]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_55_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[54]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[55]),
     .dataout(dataout[55]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_54_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[53]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[54]),
     .dataout(dataout[54]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_53_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[53]),
     .dataout(dataout[53]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_52_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[52]),
     .dataout(dataout[52]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_51_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[51]),
     .dataout(dataout[51]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_50_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[50]),
     .dataout(dataout[50]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_49_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[49]),
     .dataout(dataout[49]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_48_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[48]),
     .dataout(dataout[48]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_31_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[31]),
     .dataout(dataout[31]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_30_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[30]),
     .dataout(dataout[30]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_29_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[29]),
     .dataout(dataout[29]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_28_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[28]),
     .dataout(dataout[28]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_27_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[27]),
     .dataout(dataout[27]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_26_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[26]),
     .dataout(dataout[26]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_25_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[25]),
     .dataout(dataout[25]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_24_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[24]),
     .dataout(dataout[24]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_23_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[23]),
     .dataout(dataout[23]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_22_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[22]),
     .dataout(dataout[22]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_21_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[21]),
     .dataout(dataout[21]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_20_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[20]),
     .dataout(dataout[20]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_19_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[19]),
     .dataout(dataout[19]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_18_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[18]),
     .dataout(dataout[18]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_17_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[17]),
     .dataout(dataout[17]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_16_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[16]),
     .dataout(dataout[16]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_powersurg_buf I161 ( .in(cram_write), .o(net104));
ml_powersurg_buf I165 ( .in(net108), .o(net106));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net108));
ml_powersurg_buf I163 ( .in(net106), .o(net110));
ml_powersurg_buf I162 ( .in(net116), .o(net112));
ml_powersurg_buf I169 ( .in(net112), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net104), .o(net116));
ml_powersurg_buf I168 ( .in(net110), .o(cram_prec_out));
inv_hvt I171 ( .A(dataout[55]), .Y(net121));
inv_hvt I172 ( .A(net121), .Y(data_out));
inv_hvt I224 ( .A(net0130), .Y(ck[14]));
inv_hvt I225 ( .A(net0129), .Y(net0130));
inv_hvt I226 ( .A(net0126), .Y(net0129));
inv_hvt I229 ( .A(latch_clock), .Y(net0122));
inv_hvt I227 ( .A(net0124), .Y(net0126));
inv_hvt I228 ( .A(net0122), .Y(net0124));
mux2_hvt I197 ( .in1(net154), .in0(dataout[4]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I185 ( .in1(data_dummy_in[2]), .in0(dataout[1]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I193 ( .in1(data_dummy_in[4]), .in0(dataout[3]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I180 ( .in1(data_dummy_in[1]), .in0(dataout[0]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I188 ( .in1(data_dummy_in[3]), .in0(dataout[2]),
     .out(data_in[3]), .sel(data_muxsel1));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_1st, View - schematic
// LAST TIME SAVED: Aug 13 13:56:25 2007
// NETLIST TIME: Aug 24 09:58:59 2009
`timescale 1ns / 1ns 

module ml_blsa_tilex2_1st ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [109:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I186 ( .A(data_muxsel), .Y(net55));
inv_hvt I187 ( .A(net55), .Y(data_muxsel_buf));
inv_hvt I190 ( .A(net61), .Y(cram_pullup_buf));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net61));
inv_hvt I198 ( .A(smc_wdic_clk), .Y(net63));
inv_hvt I199 ( .A(net63), .Y(smc_wdic_clk_buf));
inv_hvt I197 ( .A(latch_clock_in), .Y(net67));
inv_hvt I196 ( .A(net67), .Y(latch_clock_out));
inv_hvt I194 ( .A(latch_reset), .Y(net71));
inv_hvt I195 ( .A(net71), .Y(latch_reset_buf));
ml_blsa_tile_1st Iml_blsa_tile_1st_0 ( .bl(bl[55:0]),
     .cram_pullup_b(cram_pullup_buf), .latch_clock(latch_clock_out),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .datain(datain), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel_buf), .cram_write(wrt_en_mid),
     .cram_prec(prec_en_mid), .data_out(data_tile),
     .cram_write_out(wrt_en_last), .cram_prec_out(prec_en_last));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blsa_tile Iml_blsa_tile_1 ( .cram_pullup_b(cram_pullup_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_wdic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[109:56]));

endmodule
// Library - xpmem, Cell - ml_blsa_bank1k, View - schematic
// LAST TIME SAVED: Jan 26 15:31:46 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ml_blsa_bank1k ( cm_sdo_u, bl, banksel, cm_sdi_u,
     cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk );


input  banksel, cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk;

output [1:0]  cm_sdo_u;

inout [331:0]  bl;

input [1:0]  cm_sdi_u;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tilex1_last Ilt_5 ( .bl(bl[331:260]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(smc_clk),
     .latch_clock_out(net142), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf), .wrt_in(net145), .prec_in(net145),
     .latch_reset(latch_reset_buf), .datain(data_out_34),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_5), .prec_out(prec_out_5),
     .data_out(cm_sdo_u[1]));
ml_blsa_tilex1 Ilt_2 ( .bl(bl[163:110]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(net179),
     .latch_clock_out(net159), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf), .wrt_in(wrt_out_34),
     .prec_in(prec_out_34), .latch_reset(latch_reset_buf),
     .datain(data_out_01), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_2),
     .prec_out(prec_out_2), .data_out(data_out_2));
ml_blsa_tilex2_bram10k Ilt_34 ( .para_en(cor_en_8bpcfg_buf),
     .para_in(sdi1_buf), .para_out(para_out), .bl(bl[259:164]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(net142),
     .latch_clock_out(net179), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret), .wrt_in(wrt_out_5),
     .prec_in(prec_out_5), .latch_reset(latch_reset_buf),
     .datain(data_out_2), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_34),
     .prec_out(prec_out_34), .data_out(data_out_34));
tiehi I267 ( .tiehi(net145));
tiehi I268 ( .tiehi(net194));
tiehi I272 ( .tiehi(net199));
tiehi I271 ( .tiehi(net195));
tiehi I273 ( .tiehi(net193));
tiehi I270 ( .tiehi(net196));
tiehi I269 ( .tiehi(net197));
ml_dff_bl I146 ( .R(latch_reset_buf), .D(para_out), .CLK(smc_clk),
     .QN(net203), .Q(net230));
nor2_hvt I254 ( .B(net205), .Y(net212), .A(cram_pullup_b));
inv_hvt I253 ( .A(cor_en_8bpcfg_b), .Y(net209));
inv_hvt I256 ( .A(banksel), .Y(net205));
inv_hvt I255 ( .A(net212), .Y(cram_pullup_logic_b));
inv_hvt I189 ( .A(smc_clk), .Y(net215));
ml_buf_ice5 I247 ( .in(cm_sdi_u[1]), .o(sdi1_buf), .sel(net199));
ml_buf_ice5 I249 ( .in(net209), .o(cor_en_8bpcfg_buf), .sel(net199));
ml_buf_ice5 I265 ( .in(net199), .o(cm_sdo_u[0]), .sel(net230));
ml_buf_ice5 I257 ( .in(smc_wdic_clk), .o(smc_wdic_clk_buf),
     .sel(banksel));
ml_buf_ice5 I203 ( .in(data_muxsel1), .o(data_muxsel1_buf),
     .sel(banksel));
ml_buf_ice5 I205 ( .in(latch_reset), .o(latch_reset_buf),
     .sel(net193));
ml_buf_ice5 I207 ( .in(cram_write), .o(cram_write_buf), .sel(banksel));
ml_buf_ice5 I208 ( .in(cram_pullup_logic_b), .o(cram_pullup_b_buf),
     .sel(cram_pullup_logic_b));
ml_buf_ice5 I201 ( .in(cram_prec), .o(cram_prec_buf), .sel(banksel));
ml_buf_ice5 I216 ( .in(net195), .o(net217), .sel(net195));
ml_buf_ice5 I245 ( .in(cm_sdi_u[0]), .o(sdi0_buf), .sel(net199));
ml_buf_ice5 I187 ( .in(smc_clk), .o(smc_clk_buf), .sel(smc_clk));
ml_buf_ice5 I188 ( .in(net215), .o(smc_clk_buf_b_ret), .sel(net215));
ml_buf_ice5 I204 ( .in(data_muxsel), .o(data_muxsel_buf),
     .sel(banksel));
ml_buf_ice5 I227 ( .in(net197), .o(net220), .sel(net197));
nor3_hvt I217 ( .B(net196), .Y(net262), .A(net196), .C(net196));
nor3_hvt I220 ( .B(net270), .Y(net266), .A(net270), .C(net270));
nor3_hvt I218 ( .B(net262), .Y(net270), .A(net262), .C(net262));
nand3_hvt I231 ( .Y(net273), .B(net277), .C(net277), .A(net277));
nand3_hvt I230 ( .Y(net277), .B(net281), .C(net281), .A(net281));
nand3_hvt I224 ( .Y(net281), .B(net194), .C(net194), .A(net194));
ml_blsa_tilex2_1st Ilt_01 ( .wrt_in(wrt_out_2), .prec_in(prec_out_2),
     .latch_reset(latch_reset_buf), .datain(sdi0_buf),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .bl(bl[109:0]),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_01),
     .prec_out(prec_out_01), .data_out(data_out_01),
     .latch_clock_in(net159), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_out(net307), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret));

endmodule
// Library - chip, Cell - CHIP_route_top1k, View - schematic
// LAST TIME SAVED: Aug  7 13:47:32 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module CHIP_route_top1k ( cm_sdo_u1, cm_sdo_u3, bl_top,
     cm_banksel_bltld3, cm_banksel_bltrd1, cm_clk_bltld3,
     cm_clk_bltrd1, .cm_prec_bltld3(cram_prec_bltld3), cm_sdi_u1d3,
     cm_sdi_u3d2, core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3,
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1) );


input  cm_clk_bltld3, cm_clk_bltrd1, cram_prec_bltld3,
     core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1;

output [1:0]  cm_sdo_u1;
output [1:0]  cm_sdo_u3;

inout [663:0]  bl_top;

input [1:0]  cm_sdi_u1d3;
input [3:3]  cm_banksel_bltrd1;
input [1:0]  cm_sdi_u3d2;
input [1:1]  cm_banksel_bltld3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_bank1k Ibltr ( .bl(bl_top[663:332]),
     .smc_wdic_clk(smc_wdis_dclk_bltrd1), .smc_clk(cm_clk_bltrd1),
     .cm_sdi_u(cm_sdi_u3d2[1:0]), .latch_reset(core_por_b_rowu3),
     .cm_sdo_u(cm_sdo_u3[1:0]), .data_muxsel1(data_muxsel1_bltrd1),
     .data_muxsel(data_muxsel_bltrd1), .cram_write(cram_write_bltrd1),
     .cram_prec(cram_prec_bltrd1),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltrd1),
     .cram_pullup_b(cram_pullup_b_bltrd1),
     .banksel(cm_banksel_bltrd1[3]));
ml_blsa_bank1k Ibltlu1 ( .bl({bl_top[0], bl_top[1], bl_top[2],
     bl_top[3], bl_top[4], bl_top[5], bl_top[6], bl_top[7], bl_top[8],
     bl_top[9], bl_top[10], bl_top[11], bl_top[12], bl_top[13],
     bl_top[14], bl_top[15], bl_top[16], bl_top[17], bl_top[18],
     bl_top[19], bl_top[20], bl_top[21], bl_top[22], bl_top[23],
     bl_top[24], bl_top[25], bl_top[26], bl_top[27], bl_top[28],
     bl_top[29], bl_top[30], bl_top[31], bl_top[32], bl_top[33],
     bl_top[34], bl_top[35], bl_top[36], bl_top[37], bl_top[38],
     bl_top[39], bl_top[40], bl_top[41], bl_top[42], bl_top[43],
     bl_top[44], bl_top[45], bl_top[46], bl_top[47], bl_top[48],
     bl_top[49], bl_top[50], bl_top[51], bl_top[52], bl_top[53],
     bl_top[54], bl_top[55], bl_top[56], bl_top[57], bl_top[58],
     bl_top[59], bl_top[60], bl_top[61], bl_top[62], bl_top[63],
     bl_top[64], bl_top[65], bl_top[66], bl_top[67], bl_top[68],
     bl_top[69], bl_top[70], bl_top[71], bl_top[72], bl_top[73],
     bl_top[74], bl_top[75], bl_top[76], bl_top[77], bl_top[78],
     bl_top[79], bl_top[80], bl_top[81], bl_top[82], bl_top[83],
     bl_top[84], bl_top[85], bl_top[86], bl_top[87], bl_top[88],
     bl_top[89], bl_top[90], bl_top[91], bl_top[92], bl_top[93],
     bl_top[94], bl_top[95], bl_top[96], bl_top[97], bl_top[98],
     bl_top[99], bl_top[100], bl_top[101], bl_top[102], bl_top[103],
     bl_top[104], bl_top[105], bl_top[106], bl_top[107], bl_top[108],
     bl_top[109], bl_top[110], bl_top[111], bl_top[112], bl_top[113],
     bl_top[114], bl_top[115], bl_top[116], bl_top[117], bl_top[118],
     bl_top[119], bl_top[120], bl_top[121], bl_top[122], bl_top[123],
     bl_top[124], bl_top[125], bl_top[126], bl_top[127], bl_top[128],
     bl_top[129], bl_top[130], bl_top[131], bl_top[132], bl_top[133],
     bl_top[134], bl_top[135], bl_top[136], bl_top[137], bl_top[138],
     bl_top[139], bl_top[140], bl_top[141], bl_top[142], bl_top[143],
     bl_top[144], bl_top[145], bl_top[146], bl_top[147], bl_top[148],
     bl_top[149], bl_top[150], bl_top[151], bl_top[152], bl_top[153],
     bl_top[154], bl_top[155], bl_top[156], bl_top[157], bl_top[158],
     bl_top[159], bl_top[160], bl_top[161], bl_top[162], bl_top[163],
     bl_top[164], bl_top[165], bl_top[166], bl_top[167], bl_top[168],
     bl_top[169], bl_top[170], bl_top[171], bl_top[172], bl_top[173],
     bl_top[174], bl_top[175], bl_top[176], bl_top[177], bl_top[178],
     bl_top[179], bl_top[180], bl_top[181], bl_top[182], bl_top[183],
     bl_top[184], bl_top[185], bl_top[186], bl_top[187], bl_top[188],
     bl_top[189], bl_top[190], bl_top[191], bl_top[192], bl_top[193],
     bl_top[194], bl_top[195], bl_top[196], bl_top[197], bl_top[198],
     bl_top[199], bl_top[200], bl_top[201], bl_top[202], bl_top[203],
     bl_top[204], bl_top[205], bl_top[206], bl_top[207], bl_top[208],
     bl_top[209], bl_top[210], bl_top[211], bl_top[212], bl_top[213],
     bl_top[214], bl_top[215], bl_top[216], bl_top[217], bl_top[218],
     bl_top[219], bl_top[220], bl_top[221], bl_top[222], bl_top[223],
     bl_top[224], bl_top[225], bl_top[226], bl_top[227], bl_top[228],
     bl_top[229], bl_top[230], bl_top[231], bl_top[232], bl_top[233],
     bl_top[234], bl_top[235], bl_top[236], bl_top[237], bl_top[238],
     bl_top[239], bl_top[240], bl_top[241], bl_top[242], bl_top[243],
     bl_top[244], bl_top[245], bl_top[246], bl_top[247], bl_top[248],
     bl_top[249], bl_top[250], bl_top[251], bl_top[252], bl_top[253],
     bl_top[254], bl_top[255], bl_top[256], bl_top[257], bl_top[258],
     bl_top[259], bl_top[260], bl_top[261], bl_top[262], bl_top[263],
     bl_top[264], bl_top[265], bl_top[266], bl_top[267], bl_top[268],
     bl_top[269], bl_top[270], bl_top[271], bl_top[272], bl_top[273],
     bl_top[274], bl_top[275], bl_top[276], bl_top[277], bl_top[278],
     bl_top[279], bl_top[280], bl_top[281], bl_top[282], bl_top[283],
     bl_top[284], bl_top[285], bl_top[286], bl_top[287], bl_top[288],
     bl_top[289], bl_top[290], bl_top[291], bl_top[292], bl_top[293],
     bl_top[294], bl_top[295], bl_top[296], bl_top[297], bl_top[298],
     bl_top[299], bl_top[300], bl_top[301], bl_top[302], bl_top[303],
     bl_top[304], bl_top[305], bl_top[306], bl_top[307], bl_top[308],
     bl_top[309], bl_top[310], bl_top[311], bl_top[312], bl_top[313],
     bl_top[314], bl_top[315], bl_top[316], bl_top[317], bl_top[318],
     bl_top[319], bl_top[320], bl_top[321], bl_top[322], bl_top[323],
     bl_top[324], bl_top[325], bl_top[326], bl_top[327], bl_top[328],
     bl_top[329], bl_top[330], bl_top[331]}),
     .smc_wdic_clk(smc_wdis_dclk_bltld3), .smc_clk(cm_clk_bltld3),
     .cm_sdi_u(cm_sdi_u1d3[1:0]), .latch_reset(core_por_b_rowu1),
     .cm_sdo_u(cm_sdo_u1[1:0]), .data_muxsel1(data_muxsel1_bltld3),
     .data_muxsel(data_muxsel_bltld3), .cram_write(cram_write_bltld3),
     .cram_prec(cram_prec_bltld3),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltld3),
     .cram_pullup_b(cram_pullup_bltld3),
     .banksel(cm_banksel_bltld3[1]));

endmodule
// Library - xpmem, Cell - sg_bufx10bot, View - schematic
// LAST TIME SAVED: Sep 18 11:01:27 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module sg_bufx10bot ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - chip, Cell - CHIP_route_bot1k, View - schematic
// LAST TIME SAVED: May 29 13:45:36 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module CHIP_route_bot1k ( cm_banksel_blbld1_0_, cm_banksel_blbld_1_,
     cm_clk_blbld, cm_sdi_u1d, cm_sdo_u0d1, cm_sdo_u1d3, cm_sdo_u2d1,
     core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, last_rsr3, monitor_celld4,
     row_testl1, smc_core_por_bottom1, smc_core_por_bottom2,
     smc_row_incl0, smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0,
     tck_padl0, bl_bot, cm_banksel, cm_banksel_blbrd_2_, cm_clk_blbrd,
     cm_sdi_u0, cm_sdi_u1, cm_sdi_u2d, cm_sdo_u1d1, core_por_b0,
     core_por_b_rowu2, core_por_bb, core_por_rowu0, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, monitor_celld2,
     row_test0, smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd,
     smc_write, vddio_botbank, vddio_spi );
output  cm_banksel_blbld1_0_, cm_banksel_blbld_1_, cm_clk_blbld,
     core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, last_rsr3, row_testl1,
     smc_core_por_bottom1, smc_core_por_bottom2, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;


input  cm_banksel_blbrd_2_, cm_clk_blbrd, core_por_b0,
     core_por_b_rowu2, core_por_bb, core_por_rowu0, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, row_test0,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     vddio_botbank, vddio_spi;

output [1:0]  cm_sdi_u1d;
output [1:0]  cm_sdo_u1d3;
output [1:0]  cm_sdo_u2d1;
output [1:0]  cm_sdo_u0d1;
output [1:0]  monitor_celld4;

inout [663:0]  bl_bot;

input [1:0]  monitor_celld2;
input [1:0]  cm_sdi_u1;
input [1:0]  cm_sdi_u0;
input [1:0]  cm_sdo_u1d1;
input [1:0]  cm_sdi_u2d;
input [1:0]  cm_banksel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net317;

wire  [1:0]  cm_sdo_u2;

wire  [1:0]  dff_u2_d1;

wire  [1:0]  monitor_celld3;

wire  [1:0]  dff_u1_d1;

wire  [1:0]  cm_sdo_u1_buf;

wire  [1:0]  cm_sdo_u0_buf;

wire  [0:1]  net234;

wire  [0:1]  net236;

wire  [1:0]  dff_u0_d1;

wire  [1:0]  cm_sdo_u0;

wire  [1:0]  dff_u0_d0;

wire  [1:0]  cm_sdi_u0d1;

wire  [2:2]  cm_banksel_blbrd1;

wire  [1:0]  dff_u2_d0;

wire  [0:1]  net341;

wire  [1:0]  cm_sdi_u2d_buf;

wire  [0:1]  net263;

wire  [0:1]  net323;

wire  [0:1]  net233;

wire  [0:1]  net235;

wire  [0:1]  net237;



ml_blsa_bank1k Iblbr ( .bl(bl_bot[663:332]),
     .smc_wdic_clk(predata_smc_wdis_dclk),
     .smc_clk(predata_smc_clk_out), .cm_sdi_u(cm_sdi_u2d_buf[1:0]),
     .latch_reset(core_por_b_rowu2), .cm_sdo_u(cm_sdo_u2[1:0]),
     .data_muxsel1(predata_muxsel1), .data_muxsel(predata_muxsel),
     .cram_write(predata_cram_write), .cram_prec(predata_cram_prec),
     .cor_en_8bpcfg_b(predata_en_8bconfig_b),
     .cram_pullup_b(predata_cram_pullup_b),
     .banksel(cm_banksel_blbrd1[2]));
ml_blsa_bank1k Iblbl ( .bl({bl_bot[0], bl_bot[1], bl_bot[2], bl_bot[3],
     bl_bot[4], bl_bot[5], bl_bot[6], bl_bot[7], bl_bot[8], bl_bot[9],
     bl_bot[10], bl_bot[11], bl_bot[12], bl_bot[13], bl_bot[14],
     bl_bot[15], bl_bot[16], bl_bot[17], bl_bot[18], bl_bot[19],
     bl_bot[20], bl_bot[21], bl_bot[22], bl_bot[23], bl_bot[24],
     bl_bot[25], bl_bot[26], bl_bot[27], bl_bot[28], bl_bot[29],
     bl_bot[30], bl_bot[31], bl_bot[32], bl_bot[33], bl_bot[34],
     bl_bot[35], bl_bot[36], bl_bot[37], bl_bot[38], bl_bot[39],
     bl_bot[40], bl_bot[41], bl_bot[42], bl_bot[43], bl_bot[44],
     bl_bot[45], bl_bot[46], bl_bot[47], bl_bot[48], bl_bot[49],
     bl_bot[50], bl_bot[51], bl_bot[52], bl_bot[53], bl_bot[54],
     bl_bot[55], bl_bot[56], bl_bot[57], bl_bot[58], bl_bot[59],
     bl_bot[60], bl_bot[61], bl_bot[62], bl_bot[63], bl_bot[64],
     bl_bot[65], bl_bot[66], bl_bot[67], bl_bot[68], bl_bot[69],
     bl_bot[70], bl_bot[71], bl_bot[72], bl_bot[73], bl_bot[74],
     bl_bot[75], bl_bot[76], bl_bot[77], bl_bot[78], bl_bot[79],
     bl_bot[80], bl_bot[81], bl_bot[82], bl_bot[83], bl_bot[84],
     bl_bot[85], bl_bot[86], bl_bot[87], bl_bot[88], bl_bot[89],
     bl_bot[90], bl_bot[91], bl_bot[92], bl_bot[93], bl_bot[94],
     bl_bot[95], bl_bot[96], bl_bot[97], bl_bot[98], bl_bot[99],
     bl_bot[100], bl_bot[101], bl_bot[102], bl_bot[103], bl_bot[104],
     bl_bot[105], bl_bot[106], bl_bot[107], bl_bot[108], bl_bot[109],
     bl_bot[110], bl_bot[111], bl_bot[112], bl_bot[113], bl_bot[114],
     bl_bot[115], bl_bot[116], bl_bot[117], bl_bot[118], bl_bot[119],
     bl_bot[120], bl_bot[121], bl_bot[122], bl_bot[123], bl_bot[124],
     bl_bot[125], bl_bot[126], bl_bot[127], bl_bot[128], bl_bot[129],
     bl_bot[130], bl_bot[131], bl_bot[132], bl_bot[133], bl_bot[134],
     bl_bot[135], bl_bot[136], bl_bot[137], bl_bot[138], bl_bot[139],
     bl_bot[140], bl_bot[141], bl_bot[142], bl_bot[143], bl_bot[144],
     bl_bot[145], bl_bot[146], bl_bot[147], bl_bot[148], bl_bot[149],
     bl_bot[150], bl_bot[151], bl_bot[152], bl_bot[153], bl_bot[154],
     bl_bot[155], bl_bot[156], bl_bot[157], bl_bot[158], bl_bot[159],
     bl_bot[160], bl_bot[161], bl_bot[162], bl_bot[163], bl_bot[164],
     bl_bot[165], bl_bot[166], bl_bot[167], bl_bot[168], bl_bot[169],
     bl_bot[170], bl_bot[171], bl_bot[172], bl_bot[173], bl_bot[174],
     bl_bot[175], bl_bot[176], bl_bot[177], bl_bot[178], bl_bot[179],
     bl_bot[180], bl_bot[181], bl_bot[182], bl_bot[183], bl_bot[184],
     bl_bot[185], bl_bot[186], bl_bot[187], bl_bot[188], bl_bot[189],
     bl_bot[190], bl_bot[191], bl_bot[192], bl_bot[193], bl_bot[194],
     bl_bot[195], bl_bot[196], bl_bot[197], bl_bot[198], bl_bot[199],
     bl_bot[200], bl_bot[201], bl_bot[202], bl_bot[203], bl_bot[204],
     bl_bot[205], bl_bot[206], bl_bot[207], bl_bot[208], bl_bot[209],
     bl_bot[210], bl_bot[211], bl_bot[212], bl_bot[213], bl_bot[214],
     bl_bot[215], bl_bot[216], bl_bot[217], bl_bot[218], bl_bot[219],
     bl_bot[220], bl_bot[221], bl_bot[222], bl_bot[223], bl_bot[224],
     bl_bot[225], bl_bot[226], bl_bot[227], bl_bot[228], bl_bot[229],
     bl_bot[230], bl_bot[231], bl_bot[232], bl_bot[233], bl_bot[234],
     bl_bot[235], bl_bot[236], bl_bot[237], bl_bot[238], bl_bot[239],
     bl_bot[240], bl_bot[241], bl_bot[242], bl_bot[243], bl_bot[244],
     bl_bot[245], bl_bot[246], bl_bot[247], bl_bot[248], bl_bot[249],
     bl_bot[250], bl_bot[251], bl_bot[252], bl_bot[253], bl_bot[254],
     bl_bot[255], bl_bot[256], bl_bot[257], bl_bot[258], bl_bot[259],
     bl_bot[260], bl_bot[261], bl_bot[262], bl_bot[263], bl_bot[264],
     bl_bot[265], bl_bot[266], bl_bot[267], bl_bot[268], bl_bot[269],
     bl_bot[270], bl_bot[271], bl_bot[272], bl_bot[273], bl_bot[274],
     bl_bot[275], bl_bot[276], bl_bot[277], bl_bot[278], bl_bot[279],
     bl_bot[280], bl_bot[281], bl_bot[282], bl_bot[283], bl_bot[284],
     bl_bot[285], bl_bot[286], bl_bot[287], bl_bot[288], bl_bot[289],
     bl_bot[290], bl_bot[291], bl_bot[292], bl_bot[293], bl_bot[294],
     bl_bot[295], bl_bot[296], bl_bot[297], bl_bot[298], bl_bot[299],
     bl_bot[300], bl_bot[301], bl_bot[302], bl_bot[303], bl_bot[304],
     bl_bot[305], bl_bot[306], bl_bot[307], bl_bot[308], bl_bot[309],
     bl_bot[310], bl_bot[311], bl_bot[312], bl_bot[313], bl_bot[314],
     bl_bot[315], bl_bot[316], bl_bot[317], bl_bot[318], bl_bot[319],
     bl_bot[320], bl_bot[321], bl_bot[322], bl_bot[323], bl_bot[324],
     bl_bot[325], bl_bot[326], bl_bot[327], bl_bot[328], bl_bot[329],
     bl_bot[330], bl_bot[331]}), .smc_wdic_clk(smc_wdis_dclk_blbld),
     .smc_clk(cm_clk_blbld), .cm_sdi_u(cm_sdi_u0d1[1:0]),
     .latch_reset(core_por_rowu0), .cm_sdo_u(cm_sdo_u0[1:0]),
     .data_muxsel1(data_muxsel1_blbld),
     .data_muxsel(data_muxsel_blbld), .cram_write(cram_write_blbld),
     .cram_prec(cram_prec_blbld),
     .cor_en_8bpcfg_b(en_8bconfig_b_blbld),
     .cram_pullup_b(cram_pullup_blbld),
     .banksel(cm_banksel_blbld1_0_));
eh_io_pup_2_new I4 ( .core_por_b(core_por_b0), .vdd_io(vddio_botbank),
     .por_b(smc_core_por_bottom1));
eh_io_pup_2_new I5 ( .core_por_b(core_por_b0), .vdd_io(vddio_spi),
     .por_b(smc_core_por_bottom2));
tielo I559_1_ ( .tielo(net233[0]));
tielo I559_0_ ( .tielo(net233[1]));
tielo I560_1_ ( .tielo(net234[0]));
tielo I560_0_ ( .tielo(net234[1]));
tielo I561_1_ ( .tielo(net235[0]));
tielo I561_0_ ( .tielo(net235[1]));
tielo I562_1_ ( .tielo(net236[0]));
tielo I562_0_ ( .tielo(net236[1]));
tielo I563_1_ ( .tielo(net237[0]));
tielo I563_0_ ( .tielo(net237[1]));
tielo I564 ( .tielo(net238));
sg_dffbuf_modified I535_1_ ( .r(net233[0]), .d(cm_sdo_u0[1]),
     .clk(net422), .dffout(dff_u0_d0[1]));
sg_dffbuf_modified I535_0_ ( .r(net233[1]), .d(cm_sdo_u0[0]),
     .clk(net422), .dffout(dff_u0_d0[0]));
sg_dffbuf_modified I546_1_ ( .r(net236[0]), .d(cm_sdo_u2[1]),
     .clk(net415), .dffout(dff_u2_d0[1]));
sg_dffbuf_modified I546_0_ ( .r(net236[1]), .d(cm_sdo_u2[0]),
     .clk(net415), .dffout(dff_u2_d0[0]));
sg_dffbuf_modified I537_1_ ( .r(net234[0]), .d(cm_sdo_u1_buf[1]),
     .clk(net412), .dffout(dff_u1_d1[1]));
sg_dffbuf_modified I537_0_ ( .r(net234[1]), .d(cm_sdo_u1_buf[0]),
     .clk(net412), .dffout(dff_u1_d1[0]));
sg_dffbuf_modified I545_1_ ( .r(net237[0]), .d(dff_u2_d0[1]),
     .clk(net416), .dffout(dff_u2_d1[1]));
sg_dffbuf_modified I545_0_ ( .r(net237[1]), .d(dff_u2_d0[0]),
     .clk(net416), .dffout(dff_u2_d1[0]));
sg_dffbuf_modified I462_1_ ( .r(net235[0]), .d(cm_sdo_u0_buf[1]),
     .clk(net412), .dffout(dff_u0_d1[1]));
sg_dffbuf_modified I462_0_ ( .r(net235[1]), .d(cm_sdo_u0_buf[0]),
     .clk(net412), .dffout(dff_u0_d1[0]));
sg_dffbuf_modified I512 ( .r(net238), .d(last_rsr2), .clk(net412),
     .dffout(net262));
sg_bufx10bot I531_1_ ( .in(net263[0]), .out(net341[0]));
sg_bufx10bot I531_0_ ( .in(net263[1]), .out(net341[1]));
sg_bufx10bot I175 ( .in(net265), .out(data_muxsel_blbld));
sg_bufx10bot I333 ( .in(j_rst_b), .out(j_rst_bl0));
sg_bufx10bot I486 ( .in(net269), .out(cram_prec_blbld));
sg_bufx10bot I492 ( .in(net271), .out(cram_write_blbld));
sg_bufx10bot I474 ( .in(net273), .out(net369));
sg_bufx10bot I496 ( .in(en_8bconfig_b_blbrd),
     .out(predata_en_8bconfig_b));
sg_bufx10bot I481 ( .in(net277), .out(cram_rstl0));
sg_bufx10bot I495 ( .in(net279), .out(en_8bconfig_b_blbld));
sg_bufx10bot I467 ( .in(predata_muxsel1), .out(net283));
sg_bufx10bot I466 ( .in(net283), .out(data_muxsel1_blbld));
sg_bufx10bot I429_1_ ( .in(monitor_celld3[1]),
     .out(monitor_celld4[1]));
sg_bufx10bot I429_0_ ( .in(monitor_celld3[0]),
     .out(monitor_celld4[0]));
sg_bufx10bot I523 ( .in(smc_clk_mid), .out(cm_clk_blbld));
sg_bufx10bot I489 ( .in(net289), .out(cram_pullup_blbld));
sg_bufx10bot I485 ( .in(cram_prec), .out(predata_cram_prec));
sg_bufx10bot I487 ( .in(predata_cram_prec), .out(net269));
sg_bufx10bot I533_1_ ( .in(cm_sdi_u1[1]), .out(net263[0]));
sg_bufx10bot I533_0_ ( .in(cm_sdi_u1[0]), .out(net263[1]));
sg_bufx10bot I527_1_ ( .in(cm_sdi_u0[1]), .out(net323[0]));
sg_bufx10bot I527_0_ ( .in(cm_sdi_u0[0]), .out(net323[1]));
sg_bufx10bot I520 ( .in(net299), .out(net343));
sg_bufx10bot I517 ( .in(net301), .out(net357));
sg_bufx10bot I493 ( .in(predata_cram_write), .out(net271));
sg_bufx10bot I505 ( .in(net305), .out(smc_rsr_rstl0));
sg_bufx10bot I509 ( .in(net307), .out(row_testl1));
sg_bufx10bot I519 ( .in(cm_banksel[0]), .out(net299));
sg_bufx10bot I491 ( .in(cram_write), .out(predata_cram_write));
sg_bufx10bot I504 ( .in(smc_rsr_rst), .out(net337));
sg_bufx10bot I494 ( .in(predata_en_8bconfig_b), .out(net279));
sg_bufx10bot I529_1_ ( .in(net317[0]), .out(cm_sdi_u0d1[1]));
sg_bufx10bot I529_0_ ( .in(net317[1]), .out(cm_sdi_u0d1[0]));
sg_bufx10bot I476 ( .in(net319), .out(cram_vddoffl0));
sg_bufx10bot I479 ( .in(cram_rst), .out(net349));
sg_bufx10bot I530_1_ ( .in(net323[0]), .out(net317[0]));
sg_bufx10bot I530_0_ ( .in(net323[1]), .out(net317[1]));
sg_bufx10bot I439 ( .in(j_tck), .out(tck_padl0));
sg_bufx10bot I510 ( .in(net327), .out(net307));
sg_bufx10bot I482 ( .in(net329), .out(cram_pgateoffl0));
sg_bufx10bot I483 ( .in(net331), .out(net329));
sg_bufx10bot I464 ( .in(predata_muxsel), .out(net265));
sg_bufx10bot I525 ( .in(cm_clk_blbrd), .out(predata_smc_clk_out));
sg_bufx10bot I503 ( .in(net337), .out(net305));
sg_bufx10bot I490 ( .in(cram_pullup_b), .out(predata_cram_pullup_b));
sg_bufx10bot I532_1_ ( .in(net341[0]), .out(cm_sdi_u1d[1]));
sg_bufx10bot I532_0_ ( .in(net341[1]), .out(cm_sdi_u1d[0]));
sg_bufx10bot I521 ( .in(net343), .out(cm_banksel_blbld1_0_));
sg_bufx10bot I465 ( .in(data_muxsel1_blbrd), .out(predata_muxsel1));
sg_bufx10bot I484 ( .in(cram_pgateoff), .out(net331));
sg_bufx10bot I480 ( .in(net349), .out(net277));
sg_bufx10bot I518 ( .in(cm_banksel[1]), .out(net301));
sg_bufx10bot I488 ( .in(predata_cram_pullup_b), .out(net289));
sg_bufx10bot I524 ( .in(predata_smc_clk_out), .out(smc_clk_mid));
sg_bufx10bot I516 ( .in(net357), .out(cm_banksel_blbld_1_));
sg_bufx10bot I470 ( .in(net359), .out(cram_wl_enl0));
sg_bufx10bot I293 ( .in(last_rsr1), .out(last_rsr2));
sg_bufx10bot I541_1_ ( .in(dff_u0_d1[1]), .out(cm_sdo_u0d1[1]));
sg_bufx10bot I541_0_ ( .in(dff_u0_d1[0]), .out(cm_sdo_u0d1[0]));
sg_bufx10bot I539_1_ ( .in(cm_sdo_u1d1[1]), .out(cm_sdo_u1_buf[1]));
sg_bufx10bot I539_0_ ( .in(cm_sdo_u1d1[0]), .out(cm_sdo_u1_buf[0]));
sg_bufx10bot I455 ( .in(data_muxsel_blbrd), .out(predata_muxsel));
sg_bufx10bot I475 ( .in(net369), .out(smc_writel0));
sg_bufx10bot I526_1_ ( .in(cm_sdi_u2d[1]), .out(cm_sdi_u2d_buf[1]));
sg_bufx10bot I526_0_ ( .in(cm_sdi_u2d[0]), .out(cm_sdi_u2d_buf[0]));
sg_bufx10bot I459 ( .in(smc_row_inc), .out(net401));
sg_bufx10bot I477 ( .in(net375), .out(net319));
sg_bufx10bot I543_1_ ( .in(dff_u0_d0[1]), .out(cm_sdo_u0_buf[1]));
sg_bufx10bot I543_0_ ( .in(dff_u0_d0[0]), .out(cm_sdo_u0_buf[0]));
sg_bufx10bot I469 ( .in(net379), .out(smc_row_incl0));
sg_bufx10bot I522 ( .in(cm_banksel_blbrd_2_),
     .out(cm_banksel_blbrd1[2]));
sg_bufx10bot I427_1_ ( .in(monitor_celld2[1]),
     .out(monitor_celld3[1]));
sg_bufx10bot I427_0_ ( .in(monitor_celld2[0]),
     .out(monitor_celld3[0]));
sg_bufx10bot I540_1_ ( .in(dff_u1_d1[1]), .out(cm_sdo_u1d3[1]));
sg_bufx10bot I540_0_ ( .in(dff_u1_d1[0]), .out(cm_sdo_u1d3[0]));
sg_bufx10bot I473 ( .in(smc_write), .out(net273));
sg_bufx10bot I542 ( .in(net262), .out(last_rsr3));
sg_bufx10bot I497 ( .in(smc_wdis_dclk_blbrd),
     .out(predata_smc_wdis_dclk));
sg_bufx10bot I511 ( .in(row_test0), .out(net327));
sg_bufx10bot I498 ( .in(net395), .out(smc_wdis_dclk_blbld));
sg_bufx10bot I471 ( .in(net397), .out(net359));
sg_bufx10bot I499 ( .in(predata_smc_wdis_dclk), .out(net395));
sg_bufx10bot I330 ( .in(net401), .out(net379));
sg_bufx10bot I478 ( .in(cram_vddoff), .out(net375));
sg_bufx10bot I336 ( .in(core_por_bb), .out(core_por_bbl0));
sg_bufx10bot I472 ( .in(cram_wl_en), .out(net397));
bram_bufferx16 I534 ( .in(smc_clk_mid), .out(net412));
bram_bufferx16 I550_1_ ( .in(dff_u2_d1[1]), .out(cm_sdo_u2d1[1]));
bram_bufferx16 I550_0_ ( .in(dff_u2_d1[0]), .out(cm_sdo_u2d1[0]));
bram_bufferx16 I549 ( .in(net415), .out(net416));
bram_bufferx16 I548 ( .in(predata_smc_clk_out), .out(net415));
bram_bufferx16 I536 ( .in(cm_clk_blbld), .out(net422));

endmodule
// Library - chip, Cell - ring_route_ice1f_july16, View - schematic
// LAST TIME SAVED: Aug  7 13:47:50 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ring_route_ice1f_july16 ( bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0, ceb0,
     en_8bconfig_b, end_of_startup, gint_hz, gsr, hiz_b0, in_bbank,
     in_lbank, in_rbank, in_tbank, j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr,
     md_spi_b, mode0, pgate_l, pgate_r, psdo, reset_l, reset_r, shift0,
     spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out_b, tdo, update0,
     vdd_cntl_l, vdd_cntl_r, wl_l, wl_r, bl_bot, bl_top, cdone,
     uio_bbank, uio_lbank, uio_rbank, uio_tbank, vpp, bm_sdo_o,
     cf_bbank, cf_lbank, cf_r_ext, cf_rbank, cf_tbank, creset_b,
     fabric_out_12_00, fabric_out_13_01, fabric_out_13_02, fromsdo,
     oen_bbank, oen_lbank, oen_rbank, oen_tbank, out_bbank, out_lbank,
     out_rbank, out_tbank, spi_ss_in_bbank, spi_ss_in_r, tck, tdi,
     tiegnd, tievdd, tms, trstb );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, ceb0, en_8bconfig_b,
     end_of_startup, gint_hz, gsr, hiz_b0, j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out_b,
     tdo, update0;

inout  cdone, vpp;

input  creset_b, fabric_out_12_00, fabric_out_13_01, fabric_out_13_02,
     fromsdo, tck, tdi, tiegnd, tievdd, tms, trstb;

output [25:0]  in_lbank;
output [287:0]  wl_r;
output [287:0]  vdd_cntl_r;
output [287:0]  vdd_cntl_l;
output [287:0]  reset_l;
output [20:0]  in_rbank;
output [3:0]  last_rsr;
output [3:0]  bm_sdi_i;
output [287:0]  reset_r;
output [287:0]  pgate_r;
output [287:0]  wl_l;
output [7:1]  psdo;
output [3:0]  bm_banksel_i;
output [23:0]  in_bbank;
output [23:0]  in_tbank;
output [7:0]  bm_sa_i;
output [287:0]  pgate_l;

inout [23:0]  uio_bbank;
inout [25:0]  uio_lbank;
inout [663:0]  bl_top;
inout [20:0]  uio_rbank;
inout [23:0]  uio_tbank;
inout [663:0]  bl_bot;

input [20:0]  oen_rbank;
input [25:0]  out_lbank;
input [7:1]  spi_ss_in_r;
input [23:0]  out_tbank;
input [23:0]  oen_tbank;
input [20:0]  cf_rbank;
input [23:0]  oen_bbank;
input [27:0]  cf_lbank;
input [3:0]  bm_sdo_o;
input [25:0]  oen_lbank;
input [1:0]  cf_r_ext;
input [20:0]  out_rbank;
input [23:0]  cf_bbank;
input [21:16]  spi_ss_in_bbank;
input [23:0]  out_bbank;
input [23:0]  cf_tbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdi_u3d;

wire  [3:3]  cm_banksel_bltrd1;

wire  [1:1]  cm_banksel_bltld3;

wire  [1:0]  cm_sdi_u0;

wire  [3:2]  monitor_celldd;

wire  [1:0]  cm_sdi_u1;

wire  [1:0]  cm_banksel;

wire  [1:0]  cm_sdi_u3d2;

wire  [1:0]  monitor_celld4;

wire  [1:0]  cm_sdi_u2d;

wire  [2:2]  cm_banksel_blbrd;

wire  [1:0]  monitor_celld2;

wire  [1:1]  cm_banksel_blbld;

wire  [0:0]  cm_banksel_blbld1;

wire  [1:0]  cm_sdo_u3;

wire  [1:0]  cm_sdo_u3dd;

wire  [1:0]  cm_sdo_u1d1;

wire  [1:0]  cm_sdi_u1d;

wire  [1:0]  cm_sdo_u1d3;

wire  [1:0]  cm_sdo_u0d1;

wire  [1:0]  cm_sdo_u2d1;

wire  [1:0]  cm_sdi_u1d3;

wire  [1:0]  cm_sdo_u1;



lefbank_1k_july16 ilefbank_f1k ( .ren(cf_lbank[25:0]),
     .oen(oen_lbank[25:0]), .out(out_lbank[25:0]),
     .pad(uio_lbank[25:0]), .in(in_lbank[25:0]));
botbank_1k_july16 Iio_botcell ( .oen(oen_bbank[23:0]),
     .out(out_bbank[23:0]), .ren(cf_bbank[23:0]),
     .pad(uio_bbank[23:0]), .in(in_bbank[23:0]), .cdone_int(cdone_in),
     .cdone_out(cdone_out), .done(cdone), .ctst_b(creset_b),
     .ctst_b_int(creset_b_int));
rgtbank_1k_july16 Iright_bank ( .ren(cf_rbank[20:0]),
     .in(in_rbank[20:0]), .out(out_rbank[20:0]), .oen(oen_rbank[20:0]),
     .pad(uio_rbank[20:0]), .tdi_int(tdi_pad), .tck_int(tck_pad),
     .tms_int(tms_pad), .tdo_int(totdopad), .tdo_en(sdo_enable),
     .trstb_int(trst_pad), .Tdo(tdo), .TRSTb(trstb), .Tdi(tdi),
     .Tms(tms), .Tck(tck));
topbank_1k_july16 Iio_topcell ( .pad(uio_tbank[23:0]),
     .in(in_tbank[23:0]), .ren(cf_tbank[23:0]), .oen(oen_tbank[23:0]),
     .out(out_tbank[23:0]), .vppin(vppin), .vpp(vpp));
nvcm_smc_fsm Invcm_smc_fsm ( .creset_b_int(creset_b_int),
     .fromsdo(fromsdo), .fabric_out_13_02(fabric_out_13_02),
     .spi_clk_out(spi_clk_out), .bm_sdo_o(bm_sdo_o[3:0]),
     .update0(update0), .cm_sdi_u2d(cm_sdi_u2d[1:0]), .vpp(vppin),
     .j_tck(j_tck), .spi_ss_out_b(spi_ss_out_b),
     .spi_sdo_oe_b(spi_sdo_oe_b), .shift0(shift0), .mode0(mode0),
     .md_spi_b(md_spi_b), .cm_sdi_u3d(cm_sdi_u3d[1:0]),
     .j_rst_b(j_rst_b), .j_tdi(j_tdi),
     .fabric_out_12_00(fabric_out_12_00),
     .fabric_out_13_01(fabric_out_13_01), .hiz_b0(hiz_b0), .gsr(gsr),
     .gint_hz(gint_hz), .end_of_startup(end_of_startup),
     .bs_en0(bs_en0), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sweb_i(bm_sweb_i), .bm_sreb_i(bm_sreb_i),
     .bm_sdi_i(bm_sdi_i[3:0]), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bm_banksel_i(bm_banksel_i[3:0]), .tiegnd(tiegnd),
     .tievdd(tievdd), .ceb0(ceb0), .cm_sdo_u2d1(cm_sdo_u2d1[1:0]),
     .cm_sdo_u1d3(cm_sdo_u1d3[1:0]), .cm_sdo_u0d1(cm_sdo_u0d1[1:0]),
     .cdone_in(cdone_in), .cm_banksel_blbrd_2_(cm_banksel_blbrd[2]),
     .cram_sdi_u0(cm_sdi_u0[1:0]),
     .cm_banksel_bltrd_3_(cm_banksel_bltrd1[3]),
     .cm_banksel_bldld(cm_banksel[1:0]), .cm_sdi_u1(cm_sdi_u1[1:0]),
     .monitor_celldd(monitor_celldd[3:2]), .core_por_b0(core_por_b0),
     .core_por_bb(core_por_bb), .cram_pgateoff(cram_pgateoff),
     .sdo_enable(sdo_enable), .totdopad(totdopad), .trst_pad(trst_pad),
     .tms_pad(tms_pad), .tdi_pad(tdi_pad), .tck_pad(tck_pad),
     .row_test0(row_test0), .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .cm_clk_blbrd(cm_clk_blbrd),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_row_inc(smc_row_inc), .smc_write(smc_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .smc_rsr_rst(smc_rsr_rst),
     .cdone_out(cdone_out), .spi_ss_in_r(spi_ss_in_r[7:1]),
     .psdo(psdo[7:1]), .spi_sdo(spi_sdo),
     .en_8bconfig_b(en_8bconfig_b), .cm_sdo_u3dd(cm_sdo_u3dd[1:0]),
     .last_rsr3(last_rsr3),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .spi_ss_in_bbankd({spi_ss_in_bbank[21], spi_ss_in_bbank[20],
     spi_ss_in_bbank[19], spi_ss_in_bbank[17], spi_ss_in_bbank[16]}),
     .cram_pullup_b(cram_pullup_b), .cram_prec(cram_prec),
     .cram_write(cram_write), .monitor_celld4(monitor_celld4[1:0]));
CHIP_route_left1f I_chip_route_left ( cm_banksel_bltld3[1],
     cm_clk_bltld3, cm_sdi_u1d3[1:0], cm_sdo_u1d1[1:0],
     core_por_b_rowu0, core_por_b_rowu1, cram_prec_bltld3,
     cram_pullup_b_bltld3, cram_write_bltld3, data_muxsel1_bltld3,
     data_muxsel_bltld3, en_8bconfig_b_bltld3,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b, last_rsr0,
     last_rsr[1:0], monitor_celld2[1:0], pgate_l[287:0],
     reset_l[287:0], smc_wdis_dclk_bltld3r, vdd_cntl_l[287:0],
     wl_l[287:0], cf_lbank[26], cf_lbank[27], cm_banksel_blbld1[0],
     cm_banksel_blbld[1], cm_clk_blbld, cm_sdi_u1d[1:0],
     cm_sdo_u1[1:0], core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0);
CHIP_route_right1f I_chip_route_right ( cm_banksel_bltrd1_3_,
     cm_clk_bltrd1, cm_sdi_u3d2[1:0], cm_sdo_u3dd[1:0],
     core_por_b_rowu2, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_write_bltrd1, data_muxsel1_bltrd1,
     data_muxsel_bltrd1, en_8bconfig_b_bltrd1,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, net380,
     last_rsr[3:2], monitor_celldd[3:2], pgate_r[287:0],
     reset_r[287:0], smc_wdis_dclk_bltrd1, vdd_cntl_r[287:0],
     wl_r[287:0], cf_r_ext[0], cf_r_ext[1], cm_banksel_blbrd[2],
     cm_banksel_bltrd1[3], cm_clk_blbrd, cm_sdi_u3d[1:0],
     cm_sdo_u3[1:0], core_por_bb, cram_pgateoff, cram_prec,
     cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en, cram_write,
     data_muxsel1_blbrd, data_muxsel_blbrd, en_8bconfig_b, j_rst_b,
     row_test0, smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd,
     smc_write, j_tck);
CHIP_route_top1k Ichip_route_top ( .core_por_b_rowu1(core_por_b_rowu1),
     .cm_sdi_u1d3(cm_sdi_u1d3[1:0]), .cm_prec_bltld3(cram_prec_bltld3),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_b_bltld3),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1),
     .cram_write_bltrd1(cram_write_bltrd1),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3r),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel1_bltld3(data_muxsel1_bltld3),
     .data_muxsel_bltld3(data_muxsel_bltld3),
     .data_muxsel1_bltrd1(data_muxsel1_bltrd1),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1),
     .bl_top(bl_top[663:0]), .cm_sdo_u1(cm_sdo_u1[1:0]),
     .cm_sdo_u3(cm_sdo_u3[1:0]),
     .cm_banksel_bltld3(cm_banksel_bltld3[1]),
     .cm_banksel_bltrd1(cm_banksel_bltrd1_3_),
     .cm_clk_bltld3(cm_clk_bltld3), .cm_clk_bltrd1(cm_clk_bltrd1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]),
     .core_por_b_rowu3(core_por_b_rowu3));
CHIP_route_bot1k Ichip_route_bot ( .bl_bot(bl_bot[663:0]),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1[0]),
     .cm_banksel_blbld_1_(cm_banksel_blbld[1]),
     .cm_clk_blbld(cm_clk_blbld), .cm_sdi_u1d(cm_sdi_u1d[1:0]),
     .cm_sdo_u0d1(cm_sdo_u0d1[1:0]), .cm_sdo_u1d3(cm_sdo_u1d3[1:0]),
     .cm_sdo_u2d1(cm_sdo_u2d1[1:0]), .core_por_bbl0(core_por_bbl0),
     .cram_pgateoffl0(cram_pgateoffl0),
     .cram_prec_blbld(cram_prec_blbld),
     .cram_pullup_blbld(cram_pullup_blbld), .cram_rstl0(cram_rstl0),
     .cram_vddoffl0(cram_vddoffl0), .cram_wl_enl0(cram_wl_enl0),
     .cram_write_blbld(cram_write_blbld),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld), .j_rst_bl0(j_rst_bl0),
     .last_rsr3(last_rsr3), .monitor_celld4(monitor_celld4[1:0]),
     .row_testl1(row_testl1),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_row_incl0(smc_row_incl0), .smc_rsr_rstl0(smc_rsr_rstl0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .smc_writel0(smc_writel0), .tck_padl0(tck_padl0),
     .cm_banksel(cm_banksel[1:0]),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd[2]),
     .cm_clk_blbrd(cm_clk_blbrd), .cm_sdi_u0(cm_sdi_u0[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdo_u1d1(cm_sdo_u1d1[1:0]), .core_por_b0(core_por_b0),
     .core_por_b_rowu2(core_por_b_rowu2), .core_por_bb(core_por_bb),
     .core_por_rowu0(core_por_b_rowu0), .cram_pgateoff(cram_pgateoff),
     .cram_prec(cram_prec), .cram_pullup_b(cram_pullup_b),
     .cram_rst(cram_rst), .cram_vddoff(cram_vddoff),
     .cram_wl_en(cram_wl_en), .cram_write(cram_write),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .en_8bconfig_b_blbrd(en_8bconfig_b), .j_rst_b(j_rst_b),
     .j_tck(j_tck), .last_rsr1(last_rsr0),
     .monitor_celld2(monitor_celld2[1:0]), .row_test0(row_test0),
     .smc_row_inc(smc_row_inc), .smc_rsr_rst(smc_rsr_rst),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd), .smc_write(smc_write),
     .vddio_botbank(vddio_bottombank), .vddio_spi(vddio_spi));

endmodule
// Library - xpmem, Cell - cram2x2, View - schematic
// LAST TIME SAVED: Jul 28 08:23:43 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module cram2x2 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [3:0]  q;
output [3:0]  q_b;

inout [1:0]  bl;

input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  r_vdd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



eh_cram_cell_4 Icram_cellb831r255 ( .q_b(q_b[1]), .q(q[1]), .wl(wl[0]),
     .bl(bl[1]), .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I20 ( .q_b(q_b[2]), .q(q[2]), .wl(wl[1]), .bl(bl[0]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));
eh_cram_cell_4 I15 ( .q_b(q_b[0]), .q(q[0]), .wl(wl[0]), .bl(bl[0]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I19 ( .q_b(q_b[3]), .q(q[3]), .wl(wl[1]), .bl(bl[1]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tiehigh, View - schematic
// LAST TIME SAVED: May  8 16:23:56 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module vdd_tiehigh ( vdd_tieh );
inout  vdd_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(vdd_tieh), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - xpmem, Cell - cram2x2x2, View - schematic
// LAST TIME SAVED: Apr 14 10:22:48 2008
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module cram2x2x2 ( q, q_b, bl, pgate_l, pgate_r, r_gnd_l, r_gnd_r,
     reset_b_l, reset_b_r, wl_l, wl_r );



output [7:0]  q_b;
output [7:0]  q;

inout [3:0]  bl;

input [1:0]  reset_b_r;
input [1:0]  pgate_l;
input [1:0]  r_gnd_r;
input [1:0]  r_gnd_l;
input [1:0]  pgate_r;
input [1:0]  wl_l;
input [1:0]  reset_b_l;
input [1:0]  wl_r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imrgt ( .bl(bl[3:2]), .q_b(q_b[7:4]), .reset(reset_b_r[1:0]),
     .q(q[7:4]), .wl(wl_r[1:0]), .r_vdd(r_gnd_r[1:0]),
     .pgate(pgate_r[1:0]));
cram2x2 Imleft ( .reset(reset_b_l[1:0]), .r_vdd(r_gnd_l[1:0]),
     .pgate(pgate_l[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl_l[1:0]));

endmodule
// Library - leafcell, Cell - ice1f_cram_row142col4, View - schematic
// LAST TIME SAVED: Apr 20 11:06:50 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ice1f_cram_row142col4 ( bl, pgate_l, pgate_r, reset_l, reset_r,
     vdd_cntl_l, vdd_cntl_r, wl_l, wl_r );


inout [3:0]  bl;

input [141:0]  wl_l;
input [141:0]  pgate_r;
input [141:0]  reset_r;
input [141:0]  vdd_cntl_r;
input [141:0]  reset_l;
input [141:0]  wl_r;
input [141:0]  vdd_cntl_l;
input [141:0]  pgate_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [141:0]  r_gnd_r;

wire  [0:567]  net29;

wire  [141:0]  r_gnd_l;

wire  [0:567]  net36;



cram2x2x2 I_cram_extra334x4_70_ ( .q(net29[0:7]),
     .reset_b_l(reset_l[141:140]), .reset_b_r(reset_r[141:140]),
     .wl_r(wl_r[141:140]), .pgate_r(pgate_r[141:140]),
     .r_gnd_r(r_gnd_r[141:140]), .r_gnd_l(r_gnd_l[141:140]),
     .q_b(net36[0:7]), .wl_l(wl_l[141:140]),
     .pgate_l(pgate_l[141:140]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_69_ ( .q(net29[8:15]),
     .reset_b_l(reset_l[139:138]), .reset_b_r(reset_r[139:138]),
     .wl_r(wl_r[139:138]), .pgate_r(pgate_r[139:138]),
     .r_gnd_r(r_gnd_r[139:138]), .r_gnd_l(r_gnd_l[139:138]),
     .q_b(net36[8:15]), .wl_l(wl_l[139:138]),
     .pgate_l(pgate_l[139:138]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_68_ ( .q(net29[16:23]),
     .reset_b_l(reset_l[137:136]), .reset_b_r(reset_r[137:136]),
     .wl_r(wl_r[137:136]), .pgate_r(pgate_r[137:136]),
     .r_gnd_r(r_gnd_r[137:136]), .r_gnd_l(r_gnd_l[137:136]),
     .q_b(net36[16:23]), .wl_l(wl_l[137:136]),
     .pgate_l(pgate_l[137:136]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_67_ ( .q(net29[24:31]),
     .reset_b_l(reset_l[135:134]), .reset_b_r(reset_r[135:134]),
     .wl_r(wl_r[135:134]), .pgate_r(pgate_r[135:134]),
     .r_gnd_r(r_gnd_r[135:134]), .r_gnd_l(r_gnd_l[135:134]),
     .q_b(net36[24:31]), .wl_l(wl_l[135:134]),
     .pgate_l(pgate_l[135:134]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_66_ ( .q(net29[32:39]),
     .reset_b_l(reset_l[133:132]), .reset_b_r(reset_r[133:132]),
     .wl_r(wl_r[133:132]), .pgate_r(pgate_r[133:132]),
     .r_gnd_r(r_gnd_r[133:132]), .r_gnd_l(r_gnd_l[133:132]),
     .q_b(net36[32:39]), .wl_l(wl_l[133:132]),
     .pgate_l(pgate_l[133:132]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_65_ ( .q(net29[40:47]),
     .reset_b_l(reset_l[131:130]), .reset_b_r(reset_r[131:130]),
     .wl_r(wl_r[131:130]), .pgate_r(pgate_r[131:130]),
     .r_gnd_r(r_gnd_r[131:130]), .r_gnd_l(r_gnd_l[131:130]),
     .q_b(net36[40:47]), .wl_l(wl_l[131:130]),
     .pgate_l(pgate_l[131:130]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_64_ ( .q(net29[48:55]),
     .reset_b_l(reset_l[129:128]), .reset_b_r(reset_r[129:128]),
     .wl_r(wl_r[129:128]), .pgate_r(pgate_r[129:128]),
     .r_gnd_r(r_gnd_r[129:128]), .r_gnd_l(r_gnd_l[129:128]),
     .q_b(net36[48:55]), .wl_l(wl_l[129:128]),
     .pgate_l(pgate_l[129:128]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_63_ ( .q(net29[56:63]),
     .reset_b_l(reset_l[127:126]), .reset_b_r(reset_r[127:126]),
     .wl_r(wl_r[127:126]), .pgate_r(pgate_r[127:126]),
     .r_gnd_r(r_gnd_r[127:126]), .r_gnd_l(r_gnd_l[127:126]),
     .q_b(net36[56:63]), .wl_l(wl_l[127:126]),
     .pgate_l(pgate_l[127:126]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_62_ ( .q(net29[64:71]),
     .reset_b_l(reset_l[125:124]), .reset_b_r(reset_r[125:124]),
     .wl_r(wl_r[125:124]), .pgate_r(pgate_r[125:124]),
     .r_gnd_r(r_gnd_r[125:124]), .r_gnd_l(r_gnd_l[125:124]),
     .q_b(net36[64:71]), .wl_l(wl_l[125:124]),
     .pgate_l(pgate_l[125:124]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_61_ ( .q(net29[72:79]),
     .reset_b_l(reset_l[123:122]), .reset_b_r(reset_r[123:122]),
     .wl_r(wl_r[123:122]), .pgate_r(pgate_r[123:122]),
     .r_gnd_r(r_gnd_r[123:122]), .r_gnd_l(r_gnd_l[123:122]),
     .q_b(net36[72:79]), .wl_l(wl_l[123:122]),
     .pgate_l(pgate_l[123:122]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_60_ ( .q(net29[80:87]),
     .reset_b_l(reset_l[121:120]), .reset_b_r(reset_r[121:120]),
     .wl_r(wl_r[121:120]), .pgate_r(pgate_r[121:120]),
     .r_gnd_r(r_gnd_r[121:120]), .r_gnd_l(r_gnd_l[121:120]),
     .q_b(net36[80:87]), .wl_l(wl_l[121:120]),
     .pgate_l(pgate_l[121:120]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_59_ ( .q(net29[88:95]),
     .reset_b_l(reset_l[119:118]), .reset_b_r(reset_r[119:118]),
     .wl_r(wl_r[119:118]), .pgate_r(pgate_r[119:118]),
     .r_gnd_r(r_gnd_r[119:118]), .r_gnd_l(r_gnd_l[119:118]),
     .q_b(net36[88:95]), .wl_l(wl_l[119:118]),
     .pgate_l(pgate_l[119:118]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_58_ ( .q(net29[96:103]),
     .reset_b_l(reset_l[117:116]), .reset_b_r(reset_r[117:116]),
     .wl_r(wl_r[117:116]), .pgate_r(pgate_r[117:116]),
     .r_gnd_r(r_gnd_r[117:116]), .r_gnd_l(r_gnd_l[117:116]),
     .q_b(net36[96:103]), .wl_l(wl_l[117:116]),
     .pgate_l(pgate_l[117:116]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_57_ ( .q(net29[104:111]),
     .reset_b_l(reset_l[115:114]), .reset_b_r(reset_r[115:114]),
     .wl_r(wl_r[115:114]), .pgate_r(pgate_r[115:114]),
     .r_gnd_r(r_gnd_r[115:114]), .r_gnd_l(r_gnd_l[115:114]),
     .q_b(net36[104:111]), .wl_l(wl_l[115:114]),
     .pgate_l(pgate_l[115:114]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_56_ ( .q(net29[112:119]),
     .reset_b_l(reset_l[113:112]), .reset_b_r(reset_r[113:112]),
     .wl_r(wl_r[113:112]), .pgate_r(pgate_r[113:112]),
     .r_gnd_r(r_gnd_r[113:112]), .r_gnd_l(r_gnd_l[113:112]),
     .q_b(net36[112:119]), .wl_l(wl_l[113:112]),
     .pgate_l(pgate_l[113:112]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_55_ ( .q(net29[120:127]),
     .reset_b_l(reset_l[111:110]), .reset_b_r(reset_r[111:110]),
     .wl_r(wl_r[111:110]), .pgate_r(pgate_r[111:110]),
     .r_gnd_r(r_gnd_r[111:110]), .r_gnd_l(r_gnd_l[111:110]),
     .q_b(net36[120:127]), .wl_l(wl_l[111:110]),
     .pgate_l(pgate_l[111:110]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_54_ ( .q(net29[128:135]),
     .reset_b_l(reset_l[109:108]), .reset_b_r(reset_r[109:108]),
     .wl_r(wl_r[109:108]), .pgate_r(pgate_r[109:108]),
     .r_gnd_r(r_gnd_r[109:108]), .r_gnd_l(r_gnd_l[109:108]),
     .q_b(net36[128:135]), .wl_l(wl_l[109:108]),
     .pgate_l(pgate_l[109:108]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_53_ ( .q(net29[136:143]),
     .reset_b_l(reset_l[107:106]), .reset_b_r(reset_r[107:106]),
     .wl_r(wl_r[107:106]), .pgate_r(pgate_r[107:106]),
     .r_gnd_r(r_gnd_r[107:106]), .r_gnd_l(r_gnd_l[107:106]),
     .q_b(net36[136:143]), .wl_l(wl_l[107:106]),
     .pgate_l(pgate_l[107:106]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_52_ ( .q(net29[144:151]),
     .reset_b_l(reset_l[105:104]), .reset_b_r(reset_r[105:104]),
     .wl_r(wl_r[105:104]), .pgate_r(pgate_r[105:104]),
     .r_gnd_r(r_gnd_r[105:104]), .r_gnd_l(r_gnd_l[105:104]),
     .q_b(net36[144:151]), .wl_l(wl_l[105:104]),
     .pgate_l(pgate_l[105:104]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_51_ ( .q(net29[152:159]),
     .reset_b_l(reset_l[103:102]), .reset_b_r(reset_r[103:102]),
     .wl_r(wl_r[103:102]), .pgate_r(pgate_r[103:102]),
     .r_gnd_r(r_gnd_r[103:102]), .r_gnd_l(r_gnd_l[103:102]),
     .q_b(net36[152:159]), .wl_l(wl_l[103:102]),
     .pgate_l(pgate_l[103:102]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_50_ ( .q(net29[160:167]),
     .reset_b_l(reset_l[101:100]), .reset_b_r(reset_r[101:100]),
     .wl_r(wl_r[101:100]), .pgate_r(pgate_r[101:100]),
     .r_gnd_r(r_gnd_r[101:100]), .r_gnd_l(r_gnd_l[101:100]),
     .q_b(net36[160:167]), .wl_l(wl_l[101:100]),
     .pgate_l(pgate_l[101:100]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_49_ ( .q(net29[168:175]),
     .reset_b_l(reset_l[99:98]), .reset_b_r(reset_r[99:98]),
     .wl_r(wl_r[99:98]), .pgate_r(pgate_r[99:98]),
     .r_gnd_r(r_gnd_r[99:98]), .r_gnd_l(r_gnd_l[99:98]),
     .q_b(net36[168:175]), .wl_l(wl_l[99:98]),
     .pgate_l(pgate_l[99:98]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_48_ ( .q(net29[176:183]),
     .reset_b_l(reset_l[97:96]), .reset_b_r(reset_r[97:96]),
     .wl_r(wl_r[97:96]), .pgate_r(pgate_r[97:96]),
     .r_gnd_r(r_gnd_r[97:96]), .r_gnd_l(r_gnd_l[97:96]),
     .q_b(net36[176:183]), .wl_l(wl_l[97:96]),
     .pgate_l(pgate_l[97:96]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_47_ ( .q(net29[184:191]),
     .reset_b_l(reset_l[95:94]), .reset_b_r(reset_r[95:94]),
     .wl_r(wl_r[95:94]), .pgate_r(pgate_r[95:94]),
     .r_gnd_r(r_gnd_r[95:94]), .r_gnd_l(r_gnd_l[95:94]),
     .q_b(net36[184:191]), .wl_l(wl_l[95:94]),
     .pgate_l(pgate_l[95:94]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_46_ ( .q(net29[192:199]),
     .reset_b_l(reset_l[93:92]), .reset_b_r(reset_r[93:92]),
     .wl_r(wl_r[93:92]), .pgate_r(pgate_r[93:92]),
     .r_gnd_r(r_gnd_r[93:92]), .r_gnd_l(r_gnd_l[93:92]),
     .q_b(net36[192:199]), .wl_l(wl_l[93:92]),
     .pgate_l(pgate_l[93:92]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_45_ ( .q(net29[200:207]),
     .reset_b_l(reset_l[91:90]), .reset_b_r(reset_r[91:90]),
     .wl_r(wl_r[91:90]), .pgate_r(pgate_r[91:90]),
     .r_gnd_r(r_gnd_r[91:90]), .r_gnd_l(r_gnd_l[91:90]),
     .q_b(net36[200:207]), .wl_l(wl_l[91:90]),
     .pgate_l(pgate_l[91:90]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_44_ ( .q(net29[208:215]),
     .reset_b_l(reset_l[89:88]), .reset_b_r(reset_r[89:88]),
     .wl_r(wl_r[89:88]), .pgate_r(pgate_r[89:88]),
     .r_gnd_r(r_gnd_r[89:88]), .r_gnd_l(r_gnd_l[89:88]),
     .q_b(net36[208:215]), .wl_l(wl_l[89:88]),
     .pgate_l(pgate_l[89:88]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_43_ ( .q(net29[216:223]),
     .reset_b_l(reset_l[87:86]), .reset_b_r(reset_r[87:86]),
     .wl_r(wl_r[87:86]), .pgate_r(pgate_r[87:86]),
     .r_gnd_r(r_gnd_r[87:86]), .r_gnd_l(r_gnd_l[87:86]),
     .q_b(net36[216:223]), .wl_l(wl_l[87:86]),
     .pgate_l(pgate_l[87:86]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_42_ ( .q(net29[224:231]),
     .reset_b_l(reset_l[85:84]), .reset_b_r(reset_r[85:84]),
     .wl_r(wl_r[85:84]), .pgate_r(pgate_r[85:84]),
     .r_gnd_r(r_gnd_r[85:84]), .r_gnd_l(r_gnd_l[85:84]),
     .q_b(net36[224:231]), .wl_l(wl_l[85:84]),
     .pgate_l(pgate_l[85:84]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_41_ ( .q(net29[232:239]),
     .reset_b_l(reset_l[83:82]), .reset_b_r(reset_r[83:82]),
     .wl_r(wl_r[83:82]), .pgate_r(pgate_r[83:82]),
     .r_gnd_r(r_gnd_r[83:82]), .r_gnd_l(r_gnd_l[83:82]),
     .q_b(net36[232:239]), .wl_l(wl_l[83:82]),
     .pgate_l(pgate_l[83:82]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_40_ ( .q(net29[240:247]),
     .reset_b_l(reset_l[81:80]), .reset_b_r(reset_r[81:80]),
     .wl_r(wl_r[81:80]), .pgate_r(pgate_r[81:80]),
     .r_gnd_r(r_gnd_r[81:80]), .r_gnd_l(r_gnd_l[81:80]),
     .q_b(net36[240:247]), .wl_l(wl_l[81:80]),
     .pgate_l(pgate_l[81:80]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_39_ ( .q(net29[248:255]),
     .reset_b_l(reset_l[79:78]), .reset_b_r(reset_r[79:78]),
     .wl_r(wl_r[79:78]), .pgate_r(pgate_r[79:78]),
     .r_gnd_r(r_gnd_r[79:78]), .r_gnd_l(r_gnd_l[79:78]),
     .q_b(net36[248:255]), .wl_l(wl_l[79:78]),
     .pgate_l(pgate_l[79:78]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_38_ ( .q(net29[256:263]),
     .reset_b_l(reset_l[77:76]), .reset_b_r(reset_r[77:76]),
     .wl_r(wl_r[77:76]), .pgate_r(pgate_r[77:76]),
     .r_gnd_r(r_gnd_r[77:76]), .r_gnd_l(r_gnd_l[77:76]),
     .q_b(net36[256:263]), .wl_l(wl_l[77:76]),
     .pgate_l(pgate_l[77:76]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_37_ ( .q(net29[264:271]),
     .reset_b_l(reset_l[75:74]), .reset_b_r(reset_r[75:74]),
     .wl_r(wl_r[75:74]), .pgate_r(pgate_r[75:74]),
     .r_gnd_r(r_gnd_r[75:74]), .r_gnd_l(r_gnd_l[75:74]),
     .q_b(net36[264:271]), .wl_l(wl_l[75:74]),
     .pgate_l(pgate_l[75:74]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_36_ ( .q(net29[272:279]),
     .reset_b_l(reset_l[73:72]), .reset_b_r(reset_r[73:72]),
     .wl_r(wl_r[73:72]), .pgate_r(pgate_r[73:72]),
     .r_gnd_r(r_gnd_r[73:72]), .r_gnd_l(r_gnd_l[73:72]),
     .q_b(net36[272:279]), .wl_l(wl_l[73:72]),
     .pgate_l(pgate_l[73:72]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_35_ ( .q(net29[280:287]),
     .reset_b_l(reset_l[71:70]), .reset_b_r(reset_r[71:70]),
     .wl_r(wl_r[71:70]), .pgate_r(pgate_r[71:70]),
     .r_gnd_r(r_gnd_r[71:70]), .r_gnd_l(r_gnd_l[71:70]),
     .q_b(net36[280:287]), .wl_l(wl_l[71:70]),
     .pgate_l(pgate_l[71:70]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_34_ ( .q(net29[288:295]),
     .reset_b_l(reset_l[69:68]), .reset_b_r(reset_r[69:68]),
     .wl_r(wl_r[69:68]), .pgate_r(pgate_r[69:68]),
     .r_gnd_r(r_gnd_r[69:68]), .r_gnd_l(r_gnd_l[69:68]),
     .q_b(net36[288:295]), .wl_l(wl_l[69:68]),
     .pgate_l(pgate_l[69:68]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_33_ ( .q(net29[296:303]),
     .reset_b_l(reset_l[67:66]), .reset_b_r(reset_r[67:66]),
     .wl_r(wl_r[67:66]), .pgate_r(pgate_r[67:66]),
     .r_gnd_r(r_gnd_r[67:66]), .r_gnd_l(r_gnd_l[67:66]),
     .q_b(net36[296:303]), .wl_l(wl_l[67:66]),
     .pgate_l(pgate_l[67:66]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_32_ ( .q(net29[304:311]),
     .reset_b_l(reset_l[65:64]), .reset_b_r(reset_r[65:64]),
     .wl_r(wl_r[65:64]), .pgate_r(pgate_r[65:64]),
     .r_gnd_r(r_gnd_r[65:64]), .r_gnd_l(r_gnd_l[65:64]),
     .q_b(net36[304:311]), .wl_l(wl_l[65:64]),
     .pgate_l(pgate_l[65:64]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_31_ ( .q(net29[312:319]),
     .reset_b_l(reset_l[63:62]), .reset_b_r(reset_r[63:62]),
     .wl_r(wl_r[63:62]), .pgate_r(pgate_r[63:62]),
     .r_gnd_r(r_gnd_r[63:62]), .r_gnd_l(r_gnd_l[63:62]),
     .q_b(net36[312:319]), .wl_l(wl_l[63:62]),
     .pgate_l(pgate_l[63:62]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_30_ ( .q(net29[320:327]),
     .reset_b_l(reset_l[61:60]), .reset_b_r(reset_r[61:60]),
     .wl_r(wl_r[61:60]), .pgate_r(pgate_r[61:60]),
     .r_gnd_r(r_gnd_r[61:60]), .r_gnd_l(r_gnd_l[61:60]),
     .q_b(net36[320:327]), .wl_l(wl_l[61:60]),
     .pgate_l(pgate_l[61:60]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_29_ ( .q(net29[328:335]),
     .reset_b_l(reset_l[59:58]), .reset_b_r(reset_r[59:58]),
     .wl_r(wl_r[59:58]), .pgate_r(pgate_r[59:58]),
     .r_gnd_r(r_gnd_r[59:58]), .r_gnd_l(r_gnd_l[59:58]),
     .q_b(net36[328:335]), .wl_l(wl_l[59:58]),
     .pgate_l(pgate_l[59:58]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_28_ ( .q(net29[336:343]),
     .reset_b_l(reset_l[57:56]), .reset_b_r(reset_r[57:56]),
     .wl_r(wl_r[57:56]), .pgate_r(pgate_r[57:56]),
     .r_gnd_r(r_gnd_r[57:56]), .r_gnd_l(r_gnd_l[57:56]),
     .q_b(net36[336:343]), .wl_l(wl_l[57:56]),
     .pgate_l(pgate_l[57:56]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_27_ ( .q(net29[344:351]),
     .reset_b_l(reset_l[55:54]), .reset_b_r(reset_r[55:54]),
     .wl_r(wl_r[55:54]), .pgate_r(pgate_r[55:54]),
     .r_gnd_r(r_gnd_r[55:54]), .r_gnd_l(r_gnd_l[55:54]),
     .q_b(net36[344:351]), .wl_l(wl_l[55:54]),
     .pgate_l(pgate_l[55:54]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_26_ ( .q(net29[352:359]),
     .reset_b_l(reset_l[53:52]), .reset_b_r(reset_r[53:52]),
     .wl_r(wl_r[53:52]), .pgate_r(pgate_r[53:52]),
     .r_gnd_r(r_gnd_r[53:52]), .r_gnd_l(r_gnd_l[53:52]),
     .q_b(net36[352:359]), .wl_l(wl_l[53:52]),
     .pgate_l(pgate_l[53:52]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_25_ ( .q(net29[360:367]),
     .reset_b_l(reset_l[51:50]), .reset_b_r(reset_r[51:50]),
     .wl_r(wl_r[51:50]), .pgate_r(pgate_r[51:50]),
     .r_gnd_r(r_gnd_r[51:50]), .r_gnd_l(r_gnd_l[51:50]),
     .q_b(net36[360:367]), .wl_l(wl_l[51:50]),
     .pgate_l(pgate_l[51:50]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_24_ ( .q(net29[368:375]),
     .reset_b_l(reset_l[49:48]), .reset_b_r(reset_r[49:48]),
     .wl_r(wl_r[49:48]), .pgate_r(pgate_r[49:48]),
     .r_gnd_r(r_gnd_r[49:48]), .r_gnd_l(r_gnd_l[49:48]),
     .q_b(net36[368:375]), .wl_l(wl_l[49:48]),
     .pgate_l(pgate_l[49:48]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_23_ ( .q(net29[376:383]),
     .reset_b_l(reset_l[47:46]), .reset_b_r(reset_r[47:46]),
     .wl_r(wl_r[47:46]), .pgate_r(pgate_r[47:46]),
     .r_gnd_r(r_gnd_r[47:46]), .r_gnd_l(r_gnd_l[47:46]),
     .q_b(net36[376:383]), .wl_l(wl_l[47:46]),
     .pgate_l(pgate_l[47:46]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_22_ ( .q(net29[384:391]),
     .reset_b_l(reset_l[45:44]), .reset_b_r(reset_r[45:44]),
     .wl_r(wl_r[45:44]), .pgate_r(pgate_r[45:44]),
     .r_gnd_r(r_gnd_r[45:44]), .r_gnd_l(r_gnd_l[45:44]),
     .q_b(net36[384:391]), .wl_l(wl_l[45:44]),
     .pgate_l(pgate_l[45:44]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_21_ ( .q(net29[392:399]),
     .reset_b_l(reset_l[43:42]), .reset_b_r(reset_r[43:42]),
     .wl_r(wl_r[43:42]), .pgate_r(pgate_r[43:42]),
     .r_gnd_r(r_gnd_r[43:42]), .r_gnd_l(r_gnd_l[43:42]),
     .q_b(net36[392:399]), .wl_l(wl_l[43:42]),
     .pgate_l(pgate_l[43:42]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_20_ ( .q(net29[400:407]),
     .reset_b_l(reset_l[41:40]), .reset_b_r(reset_r[41:40]),
     .wl_r(wl_r[41:40]), .pgate_r(pgate_r[41:40]),
     .r_gnd_r(r_gnd_r[41:40]), .r_gnd_l(r_gnd_l[41:40]),
     .q_b(net36[400:407]), .wl_l(wl_l[41:40]),
     .pgate_l(pgate_l[41:40]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_19_ ( .q(net29[408:415]),
     .reset_b_l(reset_l[39:38]), .reset_b_r(reset_r[39:38]),
     .wl_r(wl_r[39:38]), .pgate_r(pgate_r[39:38]),
     .r_gnd_r(r_gnd_r[39:38]), .r_gnd_l(r_gnd_l[39:38]),
     .q_b(net36[408:415]), .wl_l(wl_l[39:38]),
     .pgate_l(pgate_l[39:38]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_18_ ( .q(net29[416:423]),
     .reset_b_l(reset_l[37:36]), .reset_b_r(reset_r[37:36]),
     .wl_r(wl_r[37:36]), .pgate_r(pgate_r[37:36]),
     .r_gnd_r(r_gnd_r[37:36]), .r_gnd_l(r_gnd_l[37:36]),
     .q_b(net36[416:423]), .wl_l(wl_l[37:36]),
     .pgate_l(pgate_l[37:36]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_17_ ( .q(net29[424:431]),
     .reset_b_l(reset_l[35:34]), .reset_b_r(reset_r[35:34]),
     .wl_r(wl_r[35:34]), .pgate_r(pgate_r[35:34]),
     .r_gnd_r(r_gnd_r[35:34]), .r_gnd_l(r_gnd_l[35:34]),
     .q_b(net36[424:431]), .wl_l(wl_l[35:34]),
     .pgate_l(pgate_l[35:34]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_16_ ( .q(net29[432:439]),
     .reset_b_l(reset_l[33:32]), .reset_b_r(reset_r[33:32]),
     .wl_r(wl_r[33:32]), .pgate_r(pgate_r[33:32]),
     .r_gnd_r(r_gnd_r[33:32]), .r_gnd_l(r_gnd_l[33:32]),
     .q_b(net36[432:439]), .wl_l(wl_l[33:32]),
     .pgate_l(pgate_l[33:32]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_15_ ( .q(net29[440:447]),
     .reset_b_l(reset_l[31:30]), .reset_b_r(reset_r[31:30]),
     .wl_r(wl_r[31:30]), .pgate_r(pgate_r[31:30]),
     .r_gnd_r(r_gnd_r[31:30]), .r_gnd_l(r_gnd_l[31:30]),
     .q_b(net36[440:447]), .wl_l(wl_l[31:30]),
     .pgate_l(pgate_l[31:30]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_14_ ( .q(net29[448:455]),
     .reset_b_l(reset_l[29:28]), .reset_b_r(reset_r[29:28]),
     .wl_r(wl_r[29:28]), .pgate_r(pgate_r[29:28]),
     .r_gnd_r(r_gnd_r[29:28]), .r_gnd_l(r_gnd_l[29:28]),
     .q_b(net36[448:455]), .wl_l(wl_l[29:28]),
     .pgate_l(pgate_l[29:28]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_13_ ( .q(net29[456:463]),
     .reset_b_l(reset_l[27:26]), .reset_b_r(reset_r[27:26]),
     .wl_r(wl_r[27:26]), .pgate_r(pgate_r[27:26]),
     .r_gnd_r(r_gnd_r[27:26]), .r_gnd_l(r_gnd_l[27:26]),
     .q_b(net36[456:463]), .wl_l(wl_l[27:26]),
     .pgate_l(pgate_l[27:26]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_12_ ( .q(net29[464:471]),
     .reset_b_l(reset_l[25:24]), .reset_b_r(reset_r[25:24]),
     .wl_r(wl_r[25:24]), .pgate_r(pgate_r[25:24]),
     .r_gnd_r(r_gnd_r[25:24]), .r_gnd_l(r_gnd_l[25:24]),
     .q_b(net36[464:471]), .wl_l(wl_l[25:24]),
     .pgate_l(pgate_l[25:24]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_11_ ( .q(net29[472:479]),
     .reset_b_l(reset_l[23:22]), .reset_b_r(reset_r[23:22]),
     .wl_r(wl_r[23:22]), .pgate_r(pgate_r[23:22]),
     .r_gnd_r(r_gnd_r[23:22]), .r_gnd_l(r_gnd_l[23:22]),
     .q_b(net36[472:479]), .wl_l(wl_l[23:22]),
     .pgate_l(pgate_l[23:22]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_10_ ( .q(net29[480:487]),
     .reset_b_l(reset_l[21:20]), .reset_b_r(reset_r[21:20]),
     .wl_r(wl_r[21:20]), .pgate_r(pgate_r[21:20]),
     .r_gnd_r(r_gnd_r[21:20]), .r_gnd_l(r_gnd_l[21:20]),
     .q_b(net36[480:487]), .wl_l(wl_l[21:20]),
     .pgate_l(pgate_l[21:20]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_9_ ( .q(net29[488:495]),
     .reset_b_l(reset_l[19:18]), .reset_b_r(reset_r[19:18]),
     .wl_r(wl_r[19:18]), .pgate_r(pgate_r[19:18]),
     .r_gnd_r(r_gnd_r[19:18]), .r_gnd_l(r_gnd_l[19:18]),
     .q_b(net36[488:495]), .wl_l(wl_l[19:18]),
     .pgate_l(pgate_l[19:18]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_8_ ( .q(net29[496:503]),
     .reset_b_l(reset_l[17:16]), .reset_b_r(reset_r[17:16]),
     .wl_r(wl_r[17:16]), .pgate_r(pgate_r[17:16]),
     .r_gnd_r(r_gnd_r[17:16]), .r_gnd_l(r_gnd_l[17:16]),
     .q_b(net36[496:503]), .wl_l(wl_l[17:16]),
     .pgate_l(pgate_l[17:16]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_7_ ( .q(net29[504:511]),
     .reset_b_l(reset_l[15:14]), .reset_b_r(reset_r[15:14]),
     .wl_r(wl_r[15:14]), .pgate_r(pgate_r[15:14]),
     .r_gnd_r(r_gnd_r[15:14]), .r_gnd_l(r_gnd_l[15:14]),
     .q_b(net36[504:511]), .wl_l(wl_l[15:14]),
     .pgate_l(pgate_l[15:14]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_6_ ( .q(net29[512:519]),
     .reset_b_l(reset_l[13:12]), .reset_b_r(reset_r[13:12]),
     .wl_r(wl_r[13:12]), .pgate_r(pgate_r[13:12]),
     .r_gnd_r(r_gnd_r[13:12]), .r_gnd_l(r_gnd_l[13:12]),
     .q_b(net36[512:519]), .wl_l(wl_l[13:12]),
     .pgate_l(pgate_l[13:12]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_5_ ( .q(net29[520:527]),
     .reset_b_l(reset_l[11:10]), .reset_b_r(reset_r[11:10]),
     .wl_r(wl_r[11:10]), .pgate_r(pgate_r[11:10]),
     .r_gnd_r(r_gnd_r[11:10]), .r_gnd_l(r_gnd_l[11:10]),
     .q_b(net36[520:527]), .wl_l(wl_l[11:10]),
     .pgate_l(pgate_l[11:10]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_4_ ( .q(net29[528:535]),
     .reset_b_l(reset_l[9:8]), .reset_b_r(reset_r[9:8]),
     .wl_r(wl_r[9:8]), .pgate_r(pgate_r[9:8]), .r_gnd_r(r_gnd_r[9:8]),
     .r_gnd_l(r_gnd_l[9:8]), .q_b(net36[528:535]), .wl_l(wl_l[9:8]),
     .pgate_l(pgate_l[9:8]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_3_ ( .q(net29[536:543]),
     .reset_b_l(reset_l[7:6]), .reset_b_r(reset_r[7:6]),
     .wl_r(wl_r[7:6]), .pgate_r(pgate_r[7:6]), .r_gnd_r(r_gnd_r[7:6]),
     .r_gnd_l(r_gnd_l[7:6]), .q_b(net36[536:543]), .wl_l(wl_l[7:6]),
     .pgate_l(pgate_l[7:6]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_2_ ( .q(net29[544:551]),
     .reset_b_l(reset_l[5:4]), .reset_b_r(reset_r[5:4]),
     .wl_r(wl_r[5:4]), .pgate_r(pgate_r[5:4]), .r_gnd_r(r_gnd_r[5:4]),
     .r_gnd_l(r_gnd_l[5:4]), .q_b(net36[544:551]), .wl_l(wl_l[5:4]),
     .pgate_l(pgate_l[5:4]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_1_ ( .q(net29[552:559]),
     .reset_b_l(reset_l[3:2]), .reset_b_r(reset_r[3:2]),
     .wl_r(wl_r[3:2]), .pgate_r(pgate_r[3:2]), .r_gnd_r(r_gnd_r[3:2]),
     .r_gnd_l(r_gnd_l[3:2]), .q_b(net36[552:559]), .wl_l(wl_l[3:2]),
     .pgate_l(pgate_l[3:2]), .bl(bl[3:0]));
cram2x2x2 I_cram_extra334x4_0_ ( .q(net29[560:567]),
     .reset_b_l(reset_l[1:0]), .reset_b_r(reset_r[1:0]),
     .wl_r(wl_r[1:0]), .pgate_r(pgate_r[1:0]), .r_gnd_r(r_gnd_r[1:0]),
     .r_gnd_l(r_gnd_l[1:0]), .q_b(net36[560:567]), .wl_l(wl_l[1:0]),
     .pgate_l(pgate_l[1:0]), .bl(bl[3:0]));
pch_hvt  M1_141_ ( .D(r_gnd_l[141]), .B(vdd_), .G(vdd_cntl_l[141]),
     .S(vdd_));
pch_hvt  M1_140_ ( .D(r_gnd_l[140]), .B(vdd_), .G(vdd_cntl_l[140]),
     .S(vdd_));
pch_hvt  M1_139_ ( .D(r_gnd_l[139]), .B(vdd_), .G(vdd_cntl_l[139]),
     .S(vdd_));
pch_hvt  M1_138_ ( .D(r_gnd_l[138]), .B(vdd_), .G(vdd_cntl_l[138]),
     .S(vdd_));
pch_hvt  M1_137_ ( .D(r_gnd_l[137]), .B(vdd_), .G(vdd_cntl_l[137]),
     .S(vdd_));
pch_hvt  M1_136_ ( .D(r_gnd_l[136]), .B(vdd_), .G(vdd_cntl_l[136]),
     .S(vdd_));
pch_hvt  M1_135_ ( .D(r_gnd_l[135]), .B(vdd_), .G(vdd_cntl_l[135]),
     .S(vdd_));
pch_hvt  M1_134_ ( .D(r_gnd_l[134]), .B(vdd_), .G(vdd_cntl_l[134]),
     .S(vdd_));
pch_hvt  M1_133_ ( .D(r_gnd_l[133]), .B(vdd_), .G(vdd_cntl_l[133]),
     .S(vdd_));
pch_hvt  M1_132_ ( .D(r_gnd_l[132]), .B(vdd_), .G(vdd_cntl_l[132]),
     .S(vdd_));
pch_hvt  M1_131_ ( .D(r_gnd_l[131]), .B(vdd_), .G(vdd_cntl_l[131]),
     .S(vdd_));
pch_hvt  M1_130_ ( .D(r_gnd_l[130]), .B(vdd_), .G(vdd_cntl_l[130]),
     .S(vdd_));
pch_hvt  M1_129_ ( .D(r_gnd_l[129]), .B(vdd_), .G(vdd_cntl_l[129]),
     .S(vdd_));
pch_hvt  M1_128_ ( .D(r_gnd_l[128]), .B(vdd_), .G(vdd_cntl_l[128]),
     .S(vdd_));
pch_hvt  M1_127_ ( .D(r_gnd_l[127]), .B(vdd_), .G(vdd_cntl_l[127]),
     .S(vdd_));
pch_hvt  M1_126_ ( .D(r_gnd_l[126]), .B(vdd_), .G(vdd_cntl_l[126]),
     .S(vdd_));
pch_hvt  M1_125_ ( .D(r_gnd_l[125]), .B(vdd_), .G(vdd_cntl_l[125]),
     .S(vdd_));
pch_hvt  M1_124_ ( .D(r_gnd_l[124]), .B(vdd_), .G(vdd_cntl_l[124]),
     .S(vdd_));
pch_hvt  M1_123_ ( .D(r_gnd_l[123]), .B(vdd_), .G(vdd_cntl_l[123]),
     .S(vdd_));
pch_hvt  M1_122_ ( .D(r_gnd_l[122]), .B(vdd_), .G(vdd_cntl_l[122]),
     .S(vdd_));
pch_hvt  M1_121_ ( .D(r_gnd_l[121]), .B(vdd_), .G(vdd_cntl_l[121]),
     .S(vdd_));
pch_hvt  M1_120_ ( .D(r_gnd_l[120]), .B(vdd_), .G(vdd_cntl_l[120]),
     .S(vdd_));
pch_hvt  M1_119_ ( .D(r_gnd_l[119]), .B(vdd_), .G(vdd_cntl_l[119]),
     .S(vdd_));
pch_hvt  M1_118_ ( .D(r_gnd_l[118]), .B(vdd_), .G(vdd_cntl_l[118]),
     .S(vdd_));
pch_hvt  M1_117_ ( .D(r_gnd_l[117]), .B(vdd_), .G(vdd_cntl_l[117]),
     .S(vdd_));
pch_hvt  M1_116_ ( .D(r_gnd_l[116]), .B(vdd_), .G(vdd_cntl_l[116]),
     .S(vdd_));
pch_hvt  M1_115_ ( .D(r_gnd_l[115]), .B(vdd_), .G(vdd_cntl_l[115]),
     .S(vdd_));
pch_hvt  M1_114_ ( .D(r_gnd_l[114]), .B(vdd_), .G(vdd_cntl_l[114]),
     .S(vdd_));
pch_hvt  M1_113_ ( .D(r_gnd_l[113]), .B(vdd_), .G(vdd_cntl_l[113]),
     .S(vdd_));
pch_hvt  M1_112_ ( .D(r_gnd_l[112]), .B(vdd_), .G(vdd_cntl_l[112]),
     .S(vdd_));
pch_hvt  M1_111_ ( .D(r_gnd_l[111]), .B(vdd_), .G(vdd_cntl_l[111]),
     .S(vdd_));
pch_hvt  M1_110_ ( .D(r_gnd_l[110]), .B(vdd_), .G(vdd_cntl_l[110]),
     .S(vdd_));
pch_hvt  M1_109_ ( .D(r_gnd_l[109]), .B(vdd_), .G(vdd_cntl_l[109]),
     .S(vdd_));
pch_hvt  M1_108_ ( .D(r_gnd_l[108]), .B(vdd_), .G(vdd_cntl_l[108]),
     .S(vdd_));
pch_hvt  M1_107_ ( .D(r_gnd_l[107]), .B(vdd_), .G(vdd_cntl_l[107]),
     .S(vdd_));
pch_hvt  M1_106_ ( .D(r_gnd_l[106]), .B(vdd_), .G(vdd_cntl_l[106]),
     .S(vdd_));
pch_hvt  M1_105_ ( .D(r_gnd_l[105]), .B(vdd_), .G(vdd_cntl_l[105]),
     .S(vdd_));
pch_hvt  M1_104_ ( .D(r_gnd_l[104]), .B(vdd_), .G(vdd_cntl_l[104]),
     .S(vdd_));
pch_hvt  M1_103_ ( .D(r_gnd_l[103]), .B(vdd_), .G(vdd_cntl_l[103]),
     .S(vdd_));
pch_hvt  M1_102_ ( .D(r_gnd_l[102]), .B(vdd_), .G(vdd_cntl_l[102]),
     .S(vdd_));
pch_hvt  M1_101_ ( .D(r_gnd_l[101]), .B(vdd_), .G(vdd_cntl_l[101]),
     .S(vdd_));
pch_hvt  M1_100_ ( .D(r_gnd_l[100]), .B(vdd_), .G(vdd_cntl_l[100]),
     .S(vdd_));
pch_hvt  M1_99_ ( .D(r_gnd_l[99]), .B(vdd_), .G(vdd_cntl_l[99]),
     .S(vdd_));
pch_hvt  M1_98_ ( .D(r_gnd_l[98]), .B(vdd_), .G(vdd_cntl_l[98]),
     .S(vdd_));
pch_hvt  M1_97_ ( .D(r_gnd_l[97]), .B(vdd_), .G(vdd_cntl_l[97]),
     .S(vdd_));
pch_hvt  M1_96_ ( .D(r_gnd_l[96]), .B(vdd_), .G(vdd_cntl_l[96]),
     .S(vdd_));
pch_hvt  M1_95_ ( .D(r_gnd_l[95]), .B(vdd_), .G(vdd_cntl_l[95]),
     .S(vdd_));
pch_hvt  M1_94_ ( .D(r_gnd_l[94]), .B(vdd_), .G(vdd_cntl_l[94]),
     .S(vdd_));
pch_hvt  M1_93_ ( .D(r_gnd_l[93]), .B(vdd_), .G(vdd_cntl_l[93]),
     .S(vdd_));
pch_hvt  M1_92_ ( .D(r_gnd_l[92]), .B(vdd_), .G(vdd_cntl_l[92]),
     .S(vdd_));
pch_hvt  M1_91_ ( .D(r_gnd_l[91]), .B(vdd_), .G(vdd_cntl_l[91]),
     .S(vdd_));
pch_hvt  M1_90_ ( .D(r_gnd_l[90]), .B(vdd_), .G(vdd_cntl_l[90]),
     .S(vdd_));
pch_hvt  M1_89_ ( .D(r_gnd_l[89]), .B(vdd_), .G(vdd_cntl_l[89]),
     .S(vdd_));
pch_hvt  M1_88_ ( .D(r_gnd_l[88]), .B(vdd_), .G(vdd_cntl_l[88]),
     .S(vdd_));
pch_hvt  M1_87_ ( .D(r_gnd_l[87]), .B(vdd_), .G(vdd_cntl_l[87]),
     .S(vdd_));
pch_hvt  M1_86_ ( .D(r_gnd_l[86]), .B(vdd_), .G(vdd_cntl_l[86]),
     .S(vdd_));
pch_hvt  M1_85_ ( .D(r_gnd_l[85]), .B(vdd_), .G(vdd_cntl_l[85]),
     .S(vdd_));
pch_hvt  M1_84_ ( .D(r_gnd_l[84]), .B(vdd_), .G(vdd_cntl_l[84]),
     .S(vdd_));
pch_hvt  M1_83_ ( .D(r_gnd_l[83]), .B(vdd_), .G(vdd_cntl_l[83]),
     .S(vdd_));
pch_hvt  M1_82_ ( .D(r_gnd_l[82]), .B(vdd_), .G(vdd_cntl_l[82]),
     .S(vdd_));
pch_hvt  M1_81_ ( .D(r_gnd_l[81]), .B(vdd_), .G(vdd_cntl_l[81]),
     .S(vdd_));
pch_hvt  M1_80_ ( .D(r_gnd_l[80]), .B(vdd_), .G(vdd_cntl_l[80]),
     .S(vdd_));
pch_hvt  M1_79_ ( .D(r_gnd_l[79]), .B(vdd_), .G(vdd_cntl_l[79]),
     .S(vdd_));
pch_hvt  M1_78_ ( .D(r_gnd_l[78]), .B(vdd_), .G(vdd_cntl_l[78]),
     .S(vdd_));
pch_hvt  M1_77_ ( .D(r_gnd_l[77]), .B(vdd_), .G(vdd_cntl_l[77]),
     .S(vdd_));
pch_hvt  M1_76_ ( .D(r_gnd_l[76]), .B(vdd_), .G(vdd_cntl_l[76]),
     .S(vdd_));
pch_hvt  M1_75_ ( .D(r_gnd_l[75]), .B(vdd_), .G(vdd_cntl_l[75]),
     .S(vdd_));
pch_hvt  M1_74_ ( .D(r_gnd_l[74]), .B(vdd_), .G(vdd_cntl_l[74]),
     .S(vdd_));
pch_hvt  M1_73_ ( .D(r_gnd_l[73]), .B(vdd_), .G(vdd_cntl_l[73]),
     .S(vdd_));
pch_hvt  M1_72_ ( .D(r_gnd_l[72]), .B(vdd_), .G(vdd_cntl_l[72]),
     .S(vdd_));
pch_hvt  M1_71_ ( .D(r_gnd_l[71]), .B(vdd_), .G(vdd_cntl_l[71]),
     .S(vdd_));
pch_hvt  M1_70_ ( .D(r_gnd_l[70]), .B(vdd_), .G(vdd_cntl_l[70]),
     .S(vdd_));
pch_hvt  M1_69_ ( .D(r_gnd_l[69]), .B(vdd_), .G(vdd_cntl_l[69]),
     .S(vdd_));
pch_hvt  M1_68_ ( .D(r_gnd_l[68]), .B(vdd_), .G(vdd_cntl_l[68]),
     .S(vdd_));
pch_hvt  M1_67_ ( .D(r_gnd_l[67]), .B(vdd_), .G(vdd_cntl_l[67]),
     .S(vdd_));
pch_hvt  M1_66_ ( .D(r_gnd_l[66]), .B(vdd_), .G(vdd_cntl_l[66]),
     .S(vdd_));
pch_hvt  M1_65_ ( .D(r_gnd_l[65]), .B(vdd_), .G(vdd_cntl_l[65]),
     .S(vdd_));
pch_hvt  M1_64_ ( .D(r_gnd_l[64]), .B(vdd_), .G(vdd_cntl_l[64]),
     .S(vdd_));
pch_hvt  M1_63_ ( .D(r_gnd_l[63]), .B(vdd_), .G(vdd_cntl_l[63]),
     .S(vdd_));
pch_hvt  M1_62_ ( .D(r_gnd_l[62]), .B(vdd_), .G(vdd_cntl_l[62]),
     .S(vdd_));
pch_hvt  M1_61_ ( .D(r_gnd_l[61]), .B(vdd_), .G(vdd_cntl_l[61]),
     .S(vdd_));
pch_hvt  M1_60_ ( .D(r_gnd_l[60]), .B(vdd_), .G(vdd_cntl_l[60]),
     .S(vdd_));
pch_hvt  M1_59_ ( .D(r_gnd_l[59]), .B(vdd_), .G(vdd_cntl_l[59]),
     .S(vdd_));
pch_hvt  M1_58_ ( .D(r_gnd_l[58]), .B(vdd_), .G(vdd_cntl_l[58]),
     .S(vdd_));
pch_hvt  M1_57_ ( .D(r_gnd_l[57]), .B(vdd_), .G(vdd_cntl_l[57]),
     .S(vdd_));
pch_hvt  M1_56_ ( .D(r_gnd_l[56]), .B(vdd_), .G(vdd_cntl_l[56]),
     .S(vdd_));
pch_hvt  M1_55_ ( .D(r_gnd_l[55]), .B(vdd_), .G(vdd_cntl_l[55]),
     .S(vdd_));
pch_hvt  M1_54_ ( .D(r_gnd_l[54]), .B(vdd_), .G(vdd_cntl_l[54]),
     .S(vdd_));
pch_hvt  M1_53_ ( .D(r_gnd_l[53]), .B(vdd_), .G(vdd_cntl_l[53]),
     .S(vdd_));
pch_hvt  M1_52_ ( .D(r_gnd_l[52]), .B(vdd_), .G(vdd_cntl_l[52]),
     .S(vdd_));
pch_hvt  M1_51_ ( .D(r_gnd_l[51]), .B(vdd_), .G(vdd_cntl_l[51]),
     .S(vdd_));
pch_hvt  M1_50_ ( .D(r_gnd_l[50]), .B(vdd_), .G(vdd_cntl_l[50]),
     .S(vdd_));
pch_hvt  M1_49_ ( .D(r_gnd_l[49]), .B(vdd_), .G(vdd_cntl_l[49]),
     .S(vdd_));
pch_hvt  M1_48_ ( .D(r_gnd_l[48]), .B(vdd_), .G(vdd_cntl_l[48]),
     .S(vdd_));
pch_hvt  M1_47_ ( .D(r_gnd_l[47]), .B(vdd_), .G(vdd_cntl_l[47]),
     .S(vdd_));
pch_hvt  M1_46_ ( .D(r_gnd_l[46]), .B(vdd_), .G(vdd_cntl_l[46]),
     .S(vdd_));
pch_hvt  M1_45_ ( .D(r_gnd_l[45]), .B(vdd_), .G(vdd_cntl_l[45]),
     .S(vdd_));
pch_hvt  M1_44_ ( .D(r_gnd_l[44]), .B(vdd_), .G(vdd_cntl_l[44]),
     .S(vdd_));
pch_hvt  M1_43_ ( .D(r_gnd_l[43]), .B(vdd_), .G(vdd_cntl_l[43]),
     .S(vdd_));
pch_hvt  M1_42_ ( .D(r_gnd_l[42]), .B(vdd_), .G(vdd_cntl_l[42]),
     .S(vdd_));
pch_hvt  M1_41_ ( .D(r_gnd_l[41]), .B(vdd_), .G(vdd_cntl_l[41]),
     .S(vdd_));
pch_hvt  M1_40_ ( .D(r_gnd_l[40]), .B(vdd_), .G(vdd_cntl_l[40]),
     .S(vdd_));
pch_hvt  M1_39_ ( .D(r_gnd_l[39]), .B(vdd_), .G(vdd_cntl_l[39]),
     .S(vdd_));
pch_hvt  M1_38_ ( .D(r_gnd_l[38]), .B(vdd_), .G(vdd_cntl_l[38]),
     .S(vdd_));
pch_hvt  M1_37_ ( .D(r_gnd_l[37]), .B(vdd_), .G(vdd_cntl_l[37]),
     .S(vdd_));
pch_hvt  M1_36_ ( .D(r_gnd_l[36]), .B(vdd_), .G(vdd_cntl_l[36]),
     .S(vdd_));
pch_hvt  M1_35_ ( .D(r_gnd_l[35]), .B(vdd_), .G(vdd_cntl_l[35]),
     .S(vdd_));
pch_hvt  M1_34_ ( .D(r_gnd_l[34]), .B(vdd_), .G(vdd_cntl_l[34]),
     .S(vdd_));
pch_hvt  M1_33_ ( .D(r_gnd_l[33]), .B(vdd_), .G(vdd_cntl_l[33]),
     .S(vdd_));
pch_hvt  M1_32_ ( .D(r_gnd_l[32]), .B(vdd_), .G(vdd_cntl_l[32]),
     .S(vdd_));
pch_hvt  M1_31_ ( .D(r_gnd_l[31]), .B(vdd_), .G(vdd_cntl_l[31]),
     .S(vdd_));
pch_hvt  M1_30_ ( .D(r_gnd_l[30]), .B(vdd_), .G(vdd_cntl_l[30]),
     .S(vdd_));
pch_hvt  M1_29_ ( .D(r_gnd_l[29]), .B(vdd_), .G(vdd_cntl_l[29]),
     .S(vdd_));
pch_hvt  M1_28_ ( .D(r_gnd_l[28]), .B(vdd_), .G(vdd_cntl_l[28]),
     .S(vdd_));
pch_hvt  M1_27_ ( .D(r_gnd_l[27]), .B(vdd_), .G(vdd_cntl_l[27]),
     .S(vdd_));
pch_hvt  M1_26_ ( .D(r_gnd_l[26]), .B(vdd_), .G(vdd_cntl_l[26]),
     .S(vdd_));
pch_hvt  M1_25_ ( .D(r_gnd_l[25]), .B(vdd_), .G(vdd_cntl_l[25]),
     .S(vdd_));
pch_hvt  M1_24_ ( .D(r_gnd_l[24]), .B(vdd_), .G(vdd_cntl_l[24]),
     .S(vdd_));
pch_hvt  M1_23_ ( .D(r_gnd_l[23]), .B(vdd_), .G(vdd_cntl_l[23]),
     .S(vdd_));
pch_hvt  M1_22_ ( .D(r_gnd_l[22]), .B(vdd_), .G(vdd_cntl_l[22]),
     .S(vdd_));
pch_hvt  M1_21_ ( .D(r_gnd_l[21]), .B(vdd_), .G(vdd_cntl_l[21]),
     .S(vdd_));
pch_hvt  M1_20_ ( .D(r_gnd_l[20]), .B(vdd_), .G(vdd_cntl_l[20]),
     .S(vdd_));
pch_hvt  M1_19_ ( .D(r_gnd_l[19]), .B(vdd_), .G(vdd_cntl_l[19]),
     .S(vdd_));
pch_hvt  M1_18_ ( .D(r_gnd_l[18]), .B(vdd_), .G(vdd_cntl_l[18]),
     .S(vdd_));
pch_hvt  M1_17_ ( .D(r_gnd_l[17]), .B(vdd_), .G(vdd_cntl_l[17]),
     .S(vdd_));
pch_hvt  M1_16_ ( .D(r_gnd_l[16]), .B(vdd_), .G(vdd_cntl_l[16]),
     .S(vdd_));
pch_hvt  M1_15_ ( .D(r_gnd_l[15]), .B(vdd_), .G(vdd_cntl_l[15]),
     .S(vdd_));
pch_hvt  M1_14_ ( .D(r_gnd_l[14]), .B(vdd_), .G(vdd_cntl_l[14]),
     .S(vdd_));
pch_hvt  M1_13_ ( .D(r_gnd_l[13]), .B(vdd_), .G(vdd_cntl_l[13]),
     .S(vdd_));
pch_hvt  M1_12_ ( .D(r_gnd_l[12]), .B(vdd_), .G(vdd_cntl_l[12]),
     .S(vdd_));
pch_hvt  M1_11_ ( .D(r_gnd_l[11]), .B(vdd_), .G(vdd_cntl_l[11]),
     .S(vdd_));
pch_hvt  M1_10_ ( .D(r_gnd_l[10]), .B(vdd_), .G(vdd_cntl_l[10]),
     .S(vdd_));
pch_hvt  M1_9_ ( .D(r_gnd_l[9]), .B(vdd_), .G(vdd_cntl_l[9]),
     .S(vdd_));
pch_hvt  M1_8_ ( .D(r_gnd_l[8]), .B(vdd_), .G(vdd_cntl_l[8]),
     .S(vdd_));
pch_hvt  M1_7_ ( .D(r_gnd_l[7]), .B(vdd_), .G(vdd_cntl_l[7]),
     .S(vdd_));
pch_hvt  M1_6_ ( .D(r_gnd_l[6]), .B(vdd_), .G(vdd_cntl_l[6]),
     .S(vdd_));
pch_hvt  M1_5_ ( .D(r_gnd_l[5]), .B(vdd_), .G(vdd_cntl_l[5]),
     .S(vdd_));
pch_hvt  M1_4_ ( .D(r_gnd_l[4]), .B(vdd_), .G(vdd_cntl_l[4]),
     .S(vdd_));
pch_hvt  M1_3_ ( .D(r_gnd_l[3]), .B(vdd_), .G(vdd_cntl_l[3]),
     .S(vdd_));
pch_hvt  M1_2_ ( .D(r_gnd_l[2]), .B(vdd_), .G(vdd_cntl_l[2]),
     .S(vdd_));
pch_hvt  M1_1_ ( .D(r_gnd_l[1]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
pch_hvt  M1_0_ ( .D(r_gnd_l[0]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));
pch_hvt  M2_141_ ( .D(r_gnd_r[141]), .B(vdd_), .G(vdd_cntl_r[141]),
     .S(vdd_));
pch_hvt  M2_140_ ( .D(r_gnd_r[140]), .B(vdd_), .G(vdd_cntl_r[140]),
     .S(vdd_));
pch_hvt  M2_139_ ( .D(r_gnd_r[139]), .B(vdd_), .G(vdd_cntl_r[139]),
     .S(vdd_));
pch_hvt  M2_138_ ( .D(r_gnd_r[138]), .B(vdd_), .G(vdd_cntl_r[138]),
     .S(vdd_));
pch_hvt  M2_137_ ( .D(r_gnd_r[137]), .B(vdd_), .G(vdd_cntl_r[137]),
     .S(vdd_));
pch_hvt  M2_136_ ( .D(r_gnd_r[136]), .B(vdd_), .G(vdd_cntl_r[136]),
     .S(vdd_));
pch_hvt  M2_135_ ( .D(r_gnd_r[135]), .B(vdd_), .G(vdd_cntl_r[135]),
     .S(vdd_));
pch_hvt  M2_134_ ( .D(r_gnd_r[134]), .B(vdd_), .G(vdd_cntl_r[134]),
     .S(vdd_));
pch_hvt  M2_133_ ( .D(r_gnd_r[133]), .B(vdd_), .G(vdd_cntl_r[133]),
     .S(vdd_));
pch_hvt  M2_132_ ( .D(r_gnd_r[132]), .B(vdd_), .G(vdd_cntl_r[132]),
     .S(vdd_));
pch_hvt  M2_131_ ( .D(r_gnd_r[131]), .B(vdd_), .G(vdd_cntl_r[131]),
     .S(vdd_));
pch_hvt  M2_130_ ( .D(r_gnd_r[130]), .B(vdd_), .G(vdd_cntl_r[130]),
     .S(vdd_));
pch_hvt  M2_129_ ( .D(r_gnd_r[129]), .B(vdd_), .G(vdd_cntl_r[129]),
     .S(vdd_));
pch_hvt  M2_128_ ( .D(r_gnd_r[128]), .B(vdd_), .G(vdd_cntl_r[128]),
     .S(vdd_));
pch_hvt  M2_127_ ( .D(r_gnd_r[127]), .B(vdd_), .G(vdd_cntl_r[127]),
     .S(vdd_));
pch_hvt  M2_126_ ( .D(r_gnd_r[126]), .B(vdd_), .G(vdd_cntl_r[126]),
     .S(vdd_));
pch_hvt  M2_125_ ( .D(r_gnd_r[125]), .B(vdd_), .G(vdd_cntl_r[125]),
     .S(vdd_));
pch_hvt  M2_124_ ( .D(r_gnd_r[124]), .B(vdd_), .G(vdd_cntl_r[124]),
     .S(vdd_));
pch_hvt  M2_123_ ( .D(r_gnd_r[123]), .B(vdd_), .G(vdd_cntl_r[123]),
     .S(vdd_));
pch_hvt  M2_122_ ( .D(r_gnd_r[122]), .B(vdd_), .G(vdd_cntl_r[122]),
     .S(vdd_));
pch_hvt  M2_121_ ( .D(r_gnd_r[121]), .B(vdd_), .G(vdd_cntl_r[121]),
     .S(vdd_));
pch_hvt  M2_120_ ( .D(r_gnd_r[120]), .B(vdd_), .G(vdd_cntl_r[120]),
     .S(vdd_));
pch_hvt  M2_119_ ( .D(r_gnd_r[119]), .B(vdd_), .G(vdd_cntl_r[119]),
     .S(vdd_));
pch_hvt  M2_118_ ( .D(r_gnd_r[118]), .B(vdd_), .G(vdd_cntl_r[118]),
     .S(vdd_));
pch_hvt  M2_117_ ( .D(r_gnd_r[117]), .B(vdd_), .G(vdd_cntl_r[117]),
     .S(vdd_));
pch_hvt  M2_116_ ( .D(r_gnd_r[116]), .B(vdd_), .G(vdd_cntl_r[116]),
     .S(vdd_));
pch_hvt  M2_115_ ( .D(r_gnd_r[115]), .B(vdd_), .G(vdd_cntl_r[115]),
     .S(vdd_));
pch_hvt  M2_114_ ( .D(r_gnd_r[114]), .B(vdd_), .G(vdd_cntl_r[114]),
     .S(vdd_));
pch_hvt  M2_113_ ( .D(r_gnd_r[113]), .B(vdd_), .G(vdd_cntl_r[113]),
     .S(vdd_));
pch_hvt  M2_112_ ( .D(r_gnd_r[112]), .B(vdd_), .G(vdd_cntl_r[112]),
     .S(vdd_));
pch_hvt  M2_111_ ( .D(r_gnd_r[111]), .B(vdd_), .G(vdd_cntl_r[111]),
     .S(vdd_));
pch_hvt  M2_110_ ( .D(r_gnd_r[110]), .B(vdd_), .G(vdd_cntl_r[110]),
     .S(vdd_));
pch_hvt  M2_109_ ( .D(r_gnd_r[109]), .B(vdd_), .G(vdd_cntl_r[109]),
     .S(vdd_));
pch_hvt  M2_108_ ( .D(r_gnd_r[108]), .B(vdd_), .G(vdd_cntl_r[108]),
     .S(vdd_));
pch_hvt  M2_107_ ( .D(r_gnd_r[107]), .B(vdd_), .G(vdd_cntl_r[107]),
     .S(vdd_));
pch_hvt  M2_106_ ( .D(r_gnd_r[106]), .B(vdd_), .G(vdd_cntl_r[106]),
     .S(vdd_));
pch_hvt  M2_105_ ( .D(r_gnd_r[105]), .B(vdd_), .G(vdd_cntl_r[105]),
     .S(vdd_));
pch_hvt  M2_104_ ( .D(r_gnd_r[104]), .B(vdd_), .G(vdd_cntl_r[104]),
     .S(vdd_));
pch_hvt  M2_103_ ( .D(r_gnd_r[103]), .B(vdd_), .G(vdd_cntl_r[103]),
     .S(vdd_));
pch_hvt  M2_102_ ( .D(r_gnd_r[102]), .B(vdd_), .G(vdd_cntl_r[102]),
     .S(vdd_));
pch_hvt  M2_101_ ( .D(r_gnd_r[101]), .B(vdd_), .G(vdd_cntl_r[101]),
     .S(vdd_));
pch_hvt  M2_100_ ( .D(r_gnd_r[100]), .B(vdd_), .G(vdd_cntl_r[100]),
     .S(vdd_));
pch_hvt  M2_99_ ( .D(r_gnd_r[99]), .B(vdd_), .G(vdd_cntl_r[99]),
     .S(vdd_));
pch_hvt  M2_98_ ( .D(r_gnd_r[98]), .B(vdd_), .G(vdd_cntl_r[98]),
     .S(vdd_));
pch_hvt  M2_97_ ( .D(r_gnd_r[97]), .B(vdd_), .G(vdd_cntl_r[97]),
     .S(vdd_));
pch_hvt  M2_96_ ( .D(r_gnd_r[96]), .B(vdd_), .G(vdd_cntl_r[96]),
     .S(vdd_));
pch_hvt  M2_95_ ( .D(r_gnd_r[95]), .B(vdd_), .G(vdd_cntl_r[95]),
     .S(vdd_));
pch_hvt  M2_94_ ( .D(r_gnd_r[94]), .B(vdd_), .G(vdd_cntl_r[94]),
     .S(vdd_));
pch_hvt  M2_93_ ( .D(r_gnd_r[93]), .B(vdd_), .G(vdd_cntl_r[93]),
     .S(vdd_));
pch_hvt  M2_92_ ( .D(r_gnd_r[92]), .B(vdd_), .G(vdd_cntl_r[92]),
     .S(vdd_));
pch_hvt  M2_91_ ( .D(r_gnd_r[91]), .B(vdd_), .G(vdd_cntl_r[91]),
     .S(vdd_));
pch_hvt  M2_90_ ( .D(r_gnd_r[90]), .B(vdd_), .G(vdd_cntl_r[90]),
     .S(vdd_));
pch_hvt  M2_89_ ( .D(r_gnd_r[89]), .B(vdd_), .G(vdd_cntl_r[89]),
     .S(vdd_));
pch_hvt  M2_88_ ( .D(r_gnd_r[88]), .B(vdd_), .G(vdd_cntl_r[88]),
     .S(vdd_));
pch_hvt  M2_87_ ( .D(r_gnd_r[87]), .B(vdd_), .G(vdd_cntl_r[87]),
     .S(vdd_));
pch_hvt  M2_86_ ( .D(r_gnd_r[86]), .B(vdd_), .G(vdd_cntl_r[86]),
     .S(vdd_));
pch_hvt  M2_85_ ( .D(r_gnd_r[85]), .B(vdd_), .G(vdd_cntl_r[85]),
     .S(vdd_));
pch_hvt  M2_84_ ( .D(r_gnd_r[84]), .B(vdd_), .G(vdd_cntl_r[84]),
     .S(vdd_));
pch_hvt  M2_83_ ( .D(r_gnd_r[83]), .B(vdd_), .G(vdd_cntl_r[83]),
     .S(vdd_));
pch_hvt  M2_82_ ( .D(r_gnd_r[82]), .B(vdd_), .G(vdd_cntl_r[82]),
     .S(vdd_));
pch_hvt  M2_81_ ( .D(r_gnd_r[81]), .B(vdd_), .G(vdd_cntl_r[81]),
     .S(vdd_));
pch_hvt  M2_80_ ( .D(r_gnd_r[80]), .B(vdd_), .G(vdd_cntl_r[80]),
     .S(vdd_));
pch_hvt  M2_79_ ( .D(r_gnd_r[79]), .B(vdd_), .G(vdd_cntl_r[79]),
     .S(vdd_));
pch_hvt  M2_78_ ( .D(r_gnd_r[78]), .B(vdd_), .G(vdd_cntl_r[78]),
     .S(vdd_));
pch_hvt  M2_77_ ( .D(r_gnd_r[77]), .B(vdd_), .G(vdd_cntl_r[77]),
     .S(vdd_));
pch_hvt  M2_76_ ( .D(r_gnd_r[76]), .B(vdd_), .G(vdd_cntl_r[76]),
     .S(vdd_));
pch_hvt  M2_75_ ( .D(r_gnd_r[75]), .B(vdd_), .G(vdd_cntl_r[75]),
     .S(vdd_));
pch_hvt  M2_74_ ( .D(r_gnd_r[74]), .B(vdd_), .G(vdd_cntl_r[74]),
     .S(vdd_));
pch_hvt  M2_73_ ( .D(r_gnd_r[73]), .B(vdd_), .G(vdd_cntl_r[73]),
     .S(vdd_));
pch_hvt  M2_72_ ( .D(r_gnd_r[72]), .B(vdd_), .G(vdd_cntl_r[72]),
     .S(vdd_));
pch_hvt  M2_71_ ( .D(r_gnd_r[71]), .B(vdd_), .G(vdd_cntl_r[71]),
     .S(vdd_));
pch_hvt  M2_70_ ( .D(r_gnd_r[70]), .B(vdd_), .G(vdd_cntl_r[70]),
     .S(vdd_));
pch_hvt  M2_69_ ( .D(r_gnd_r[69]), .B(vdd_), .G(vdd_cntl_r[69]),
     .S(vdd_));
pch_hvt  M2_68_ ( .D(r_gnd_r[68]), .B(vdd_), .G(vdd_cntl_r[68]),
     .S(vdd_));
pch_hvt  M2_67_ ( .D(r_gnd_r[67]), .B(vdd_), .G(vdd_cntl_r[67]),
     .S(vdd_));
pch_hvt  M2_66_ ( .D(r_gnd_r[66]), .B(vdd_), .G(vdd_cntl_r[66]),
     .S(vdd_));
pch_hvt  M2_65_ ( .D(r_gnd_r[65]), .B(vdd_), .G(vdd_cntl_r[65]),
     .S(vdd_));
pch_hvt  M2_64_ ( .D(r_gnd_r[64]), .B(vdd_), .G(vdd_cntl_r[64]),
     .S(vdd_));
pch_hvt  M2_63_ ( .D(r_gnd_r[63]), .B(vdd_), .G(vdd_cntl_r[63]),
     .S(vdd_));
pch_hvt  M2_62_ ( .D(r_gnd_r[62]), .B(vdd_), .G(vdd_cntl_r[62]),
     .S(vdd_));
pch_hvt  M2_61_ ( .D(r_gnd_r[61]), .B(vdd_), .G(vdd_cntl_r[61]),
     .S(vdd_));
pch_hvt  M2_60_ ( .D(r_gnd_r[60]), .B(vdd_), .G(vdd_cntl_r[60]),
     .S(vdd_));
pch_hvt  M2_59_ ( .D(r_gnd_r[59]), .B(vdd_), .G(vdd_cntl_r[59]),
     .S(vdd_));
pch_hvt  M2_58_ ( .D(r_gnd_r[58]), .B(vdd_), .G(vdd_cntl_r[58]),
     .S(vdd_));
pch_hvt  M2_57_ ( .D(r_gnd_r[57]), .B(vdd_), .G(vdd_cntl_r[57]),
     .S(vdd_));
pch_hvt  M2_56_ ( .D(r_gnd_r[56]), .B(vdd_), .G(vdd_cntl_r[56]),
     .S(vdd_));
pch_hvt  M2_55_ ( .D(r_gnd_r[55]), .B(vdd_), .G(vdd_cntl_r[55]),
     .S(vdd_));
pch_hvt  M2_54_ ( .D(r_gnd_r[54]), .B(vdd_), .G(vdd_cntl_r[54]),
     .S(vdd_));
pch_hvt  M2_53_ ( .D(r_gnd_r[53]), .B(vdd_), .G(vdd_cntl_r[53]),
     .S(vdd_));
pch_hvt  M2_52_ ( .D(r_gnd_r[52]), .B(vdd_), .G(vdd_cntl_r[52]),
     .S(vdd_));
pch_hvt  M2_51_ ( .D(r_gnd_r[51]), .B(vdd_), .G(vdd_cntl_r[51]),
     .S(vdd_));
pch_hvt  M2_50_ ( .D(r_gnd_r[50]), .B(vdd_), .G(vdd_cntl_r[50]),
     .S(vdd_));
pch_hvt  M2_49_ ( .D(r_gnd_r[49]), .B(vdd_), .G(vdd_cntl_r[49]),
     .S(vdd_));
pch_hvt  M2_48_ ( .D(r_gnd_r[48]), .B(vdd_), .G(vdd_cntl_r[48]),
     .S(vdd_));
pch_hvt  M2_47_ ( .D(r_gnd_r[47]), .B(vdd_), .G(vdd_cntl_r[47]),
     .S(vdd_));
pch_hvt  M2_46_ ( .D(r_gnd_r[46]), .B(vdd_), .G(vdd_cntl_r[46]),
     .S(vdd_));
pch_hvt  M2_45_ ( .D(r_gnd_r[45]), .B(vdd_), .G(vdd_cntl_r[45]),
     .S(vdd_));
pch_hvt  M2_44_ ( .D(r_gnd_r[44]), .B(vdd_), .G(vdd_cntl_r[44]),
     .S(vdd_));
pch_hvt  M2_43_ ( .D(r_gnd_r[43]), .B(vdd_), .G(vdd_cntl_r[43]),
     .S(vdd_));
pch_hvt  M2_42_ ( .D(r_gnd_r[42]), .B(vdd_), .G(vdd_cntl_r[42]),
     .S(vdd_));
pch_hvt  M2_41_ ( .D(r_gnd_r[41]), .B(vdd_), .G(vdd_cntl_r[41]),
     .S(vdd_));
pch_hvt  M2_40_ ( .D(r_gnd_r[40]), .B(vdd_), .G(vdd_cntl_r[40]),
     .S(vdd_));
pch_hvt  M2_39_ ( .D(r_gnd_r[39]), .B(vdd_), .G(vdd_cntl_r[39]),
     .S(vdd_));
pch_hvt  M2_38_ ( .D(r_gnd_r[38]), .B(vdd_), .G(vdd_cntl_r[38]),
     .S(vdd_));
pch_hvt  M2_37_ ( .D(r_gnd_r[37]), .B(vdd_), .G(vdd_cntl_r[37]),
     .S(vdd_));
pch_hvt  M2_36_ ( .D(r_gnd_r[36]), .B(vdd_), .G(vdd_cntl_r[36]),
     .S(vdd_));
pch_hvt  M2_35_ ( .D(r_gnd_r[35]), .B(vdd_), .G(vdd_cntl_r[35]),
     .S(vdd_));
pch_hvt  M2_34_ ( .D(r_gnd_r[34]), .B(vdd_), .G(vdd_cntl_r[34]),
     .S(vdd_));
pch_hvt  M2_33_ ( .D(r_gnd_r[33]), .B(vdd_), .G(vdd_cntl_r[33]),
     .S(vdd_));
pch_hvt  M2_32_ ( .D(r_gnd_r[32]), .B(vdd_), .G(vdd_cntl_r[32]),
     .S(vdd_));
pch_hvt  M2_31_ ( .D(r_gnd_r[31]), .B(vdd_), .G(vdd_cntl_r[31]),
     .S(vdd_));
pch_hvt  M2_30_ ( .D(r_gnd_r[30]), .B(vdd_), .G(vdd_cntl_r[30]),
     .S(vdd_));
pch_hvt  M2_29_ ( .D(r_gnd_r[29]), .B(vdd_), .G(vdd_cntl_r[29]),
     .S(vdd_));
pch_hvt  M2_28_ ( .D(r_gnd_r[28]), .B(vdd_), .G(vdd_cntl_r[28]),
     .S(vdd_));
pch_hvt  M2_27_ ( .D(r_gnd_r[27]), .B(vdd_), .G(vdd_cntl_r[27]),
     .S(vdd_));
pch_hvt  M2_26_ ( .D(r_gnd_r[26]), .B(vdd_), .G(vdd_cntl_r[26]),
     .S(vdd_));
pch_hvt  M2_25_ ( .D(r_gnd_r[25]), .B(vdd_), .G(vdd_cntl_r[25]),
     .S(vdd_));
pch_hvt  M2_24_ ( .D(r_gnd_r[24]), .B(vdd_), .G(vdd_cntl_r[24]),
     .S(vdd_));
pch_hvt  M2_23_ ( .D(r_gnd_r[23]), .B(vdd_), .G(vdd_cntl_r[23]),
     .S(vdd_));
pch_hvt  M2_22_ ( .D(r_gnd_r[22]), .B(vdd_), .G(vdd_cntl_r[22]),
     .S(vdd_));
pch_hvt  M2_21_ ( .D(r_gnd_r[21]), .B(vdd_), .G(vdd_cntl_r[21]),
     .S(vdd_));
pch_hvt  M2_20_ ( .D(r_gnd_r[20]), .B(vdd_), .G(vdd_cntl_r[20]),
     .S(vdd_));
pch_hvt  M2_19_ ( .D(r_gnd_r[19]), .B(vdd_), .G(vdd_cntl_r[19]),
     .S(vdd_));
pch_hvt  M2_18_ ( .D(r_gnd_r[18]), .B(vdd_), .G(vdd_cntl_r[18]),
     .S(vdd_));
pch_hvt  M2_17_ ( .D(r_gnd_r[17]), .B(vdd_), .G(vdd_cntl_r[17]),
     .S(vdd_));
pch_hvt  M2_16_ ( .D(r_gnd_r[16]), .B(vdd_), .G(vdd_cntl_r[16]),
     .S(vdd_));
pch_hvt  M2_15_ ( .D(r_gnd_r[15]), .B(vdd_), .G(vdd_cntl_r[15]),
     .S(vdd_));
pch_hvt  M2_14_ ( .D(r_gnd_r[14]), .B(vdd_), .G(vdd_cntl_r[14]),
     .S(vdd_));
pch_hvt  M2_13_ ( .D(r_gnd_r[13]), .B(vdd_), .G(vdd_cntl_r[13]),
     .S(vdd_));
pch_hvt  M2_12_ ( .D(r_gnd_r[12]), .B(vdd_), .G(vdd_cntl_r[12]),
     .S(vdd_));
pch_hvt  M2_11_ ( .D(r_gnd_r[11]), .B(vdd_), .G(vdd_cntl_r[11]),
     .S(vdd_));
pch_hvt  M2_10_ ( .D(r_gnd_r[10]), .B(vdd_), .G(vdd_cntl_r[10]),
     .S(vdd_));
pch_hvt  M2_9_ ( .D(r_gnd_r[9]), .B(vdd_), .G(vdd_cntl_r[9]),
     .S(vdd_));
pch_hvt  M2_8_ ( .D(r_gnd_r[8]), .B(vdd_), .G(vdd_cntl_r[8]),
     .S(vdd_));
pch_hvt  M2_7_ ( .D(r_gnd_r[7]), .B(vdd_), .G(vdd_cntl_r[7]),
     .S(vdd_));
pch_hvt  M2_6_ ( .D(r_gnd_r[6]), .B(vdd_), .G(vdd_cntl_r[6]),
     .S(vdd_));
pch_hvt  M2_5_ ( .D(r_gnd_r[5]), .B(vdd_), .G(vdd_cntl_r[5]),
     .S(vdd_));
pch_hvt  M2_4_ ( .D(r_gnd_r[4]), .B(vdd_), .G(vdd_cntl_r[4]),
     .S(vdd_));
pch_hvt  M2_3_ ( .D(r_gnd_r[3]), .B(vdd_), .G(vdd_cntl_r[3]),
     .S(vdd_));
pch_hvt  M2_2_ ( .D(r_gnd_r[2]), .B(vdd_), .G(vdd_cntl_r[2]),
     .S(vdd_));
pch_hvt  M2_1_ ( .D(r_gnd_r[1]), .B(vdd_), .G(vdd_cntl_r[1]),
     .S(vdd_));
pch_hvt  M2_0_ ( .D(r_gnd_r[0]), .B(vdd_), .G(vdd_cntl_r[0]),
     .S(vdd_));

endmodule
// Library - io, Cell - insel1_hvt_v2, View - schematic
// LAST TIME SAVED: Jul 10 10:25:59 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module insel1_hvt_v2 ( out, in0, in1, in2, in3, sb, sel );
output  out;

input  in0, in1, in2, in3;

input [1:0]  sel;
input [1:0]  sb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I39 ( .in(in3), .out(outd23), .pp(sb[0]), .nn(sel[0]));
txgate_hvt I40 ( .in(in2), .out(outd23), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I33 ( .in(outd01), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_hvt I_txgate1 ( .in(in1), .out(outd01), .pp(sb[0]),
     .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(outd01), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(outd23), .out(out), .pp(sb[1]), .nn(sel[1]));

endmodule
// Library - io, Cell - cebdffrqn, View - schematic
// LAST TIME SAVED: Jan 31 09:00:47 2008
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module cebdffrqn ( q, qn, ceb, clk, d, r );
output  q, qn;

input  ceb, clk, d, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I54 ( .A(net62), .B(clk), .Y(clatb), .C(ceb));
nand2_hvt I290 ( .A(clk), .Y(clkb), .B(clatb));
nand2_hvt I42 ( .A(si), .B(rstb), .Y(so));
nor2_hvt INAND2_m ( .A(r), .Y(q), .B(mi));
inv_hvt I39 ( .A(q), .Y(qn));
inv_hvt Iinv_ckfb ( .A(clatb), .Y(net62));
inv_hvt I50 ( .A(clkb), .Y(clkd));
inv_hvt I43 ( .A(so), .Y(low_s));
inv_hvt I40 ( .A(r), .Y(rstb));
txgate_hvt I44 ( .in(d), .out(si), .pp(clkd), .nn(clkb));
txgate_hvt I52 ( .in(so), .out(mi), .pp(clkb), .nn(clkd));
txgate_hvt I51 ( .in(si), .out(low_s), .pp(clkb), .nn(clkd));
txgate_hvt I53 ( .in(mi), .out(qn), .pp(clkd), .nn(clkb));

endmodule
// Library - io, Cell - dffrckb, View - schematic
// LAST TIME SAVED: May 11 14:58:52 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module dffrckb ( q, qn, clk, d, e, r );
output  q, qn;

input  clk, d, e, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



oai21x2_hvt I57 ( .A1(clk), .Y(clat), .A0(clatb), .B0(e));
nor2_hvt I48 ( .B(clat), .A(clk), .Y(clkb));
nand2_hvt I54 ( .A(rstb), .Y(qn), .B(q));
nand2_hvt I42 ( .A(si), .B(rstb), .Y(so));
inv_hvt I55 ( .A(mi), .Y(q));
inv_hvt I50 ( .A(clkb), .Y(clkd));
inv_hvt I56 ( .A(clat), .Y(clatb));
inv_hvt I43 ( .A(so), .Y(low_s));
inv_hvt I40 ( .A(r), .Y(rstb));
txgate_hvt I59 ( .in(d), .out(si), .pp(clkb), .nn(clkd));
txgate_hvt I64 ( .in(low_s), .out(si), .pp(clkd), .nn(clkb));
txgate_hvt I62 ( .in(qn), .out(mi), .pp(clkb), .nn(clkd));
txgate_hvt I60 ( .in(so), .out(mi), .pp(clkd), .nn(clkb));

endmodule
// Library - io, Cell - in_logic_v1rev2, View - schematic
// LAST TIME SAVED: Jul 10 10:31:59 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module in_logic_v1rev2 ( dout0, dout1, sdo, bs_en, cbit, cbitb, ceb,
     clk, cntl, din, mode, rstio, sdi, shift, tclk, ud );
output  dout0, dout1, sdo;

input  bs_en, ceb, clk, cntl, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I_inv_dout0 ( .A(doutb), .Y(dout0));
inv_hvt I_inv_dout1 ( .A(udd), .Y(dout1));
inv_hvt I185 ( .A(cbit1b), .Y(cbit1));
inv_hvt I186 ( .A(dout0), .Y(net037));
inv_hvt I172 ( .A(din), .Y(dinb));
nand2_hvt I188 ( .A(cntl), .Y(cbit1b), .B(cbit[1]));
insel1_hvt_v2 I_insel1 ( .in1(dinb), .in0(regb), .out(reg_),
     .sb({cbit1b, cbitb[0]}), .sel({cbit1, cbit[0]}), .in2(net037),
     .in3(net037));
mux2x1_hvt I_mux_mode ( .sel(mode), .in1(udd), .in0(reg_),
     .out(doutb));
cebdffrqn I_dff0 ( .ceb(ceb), .clk(ck2r0), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_dff1 ( .e(ud), .clk(ck2r0), .qn(udd), .r(rstio), .q(net060),
     .d(net056));
mux2x1_hvt I_mux_clk ( .in1(tclk), .in0(clk), .out(ck2r0),
     .sel(bs_en));
mux2x1_hvt I_mux_data ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
mux2x1_hvt I_mux2_btw ( .in1(sdo), .in0(din), .out(net056),
     .sel(bs_en));

endmodule
// Library - io, Cell - in_logic_v3rev, View - schematic
// LAST TIME SAVED: Jul 10 10:30:27 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module in_logic_v3rev ( dout0, dout1, sdo, sp12, bl, bs_en, ceb, clk,
     cntl, din, mode, pgate, prog, reset, rstio, sdi, shift, slfop,
     tclk, ud, vdd_cntl, wl );
output  dout0, dout1, sdo, sp12;


input  bs_en, ceb, clk, cntl, din, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  reset;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbit;

wire  [3:0]  cbitb;



in_logic_v1rev2 I_in_logic ( .ceb(ceb), .rstio(rstio), .din(din),
     .cntl(cntl), .dout1(dout1), .dout0(dout0), .shift(shift), .ud(ud),
     .clk(clk), .sdo(sdo), .sdi(sdi), .cbit({cbit[0], cbit[1]}),
     .cbitb({cbitb[0], cbitb[1]}), .tclk(tclk), .bs_en(bs_en),
     .mode(mode));
pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[3]), .sp12(sp12),
     .prog(prog));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - odrv12x3, View - schematic
// LAST TIME SAVED: Aug 23 11:52:00 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module odrv12x3 ( sp12, bl, pgate, prog, reset, slfop, vdd_cntl, wl );


input  prog;

output [2:0]  sp12;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  reset;
input [1:0]  vdd_cntl;
input [2:0]  slfop;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12_2_ ( .slfop(slfop[2]), .cbitb(cbitb[2]),
     .sp12(sp12[2]), .prog(prog));
odrv12 I_odrv12_1_ ( .slfop(slfop[1]), .cbitb(cbitb[1]),
     .sp12(sp12[1]), .prog(prog));
odrv12 I_odrv12_0_ ( .slfop(slfop[0]), .cbitb(cbitb[0]),
     .sp12(sp12[0]), .prog(prog));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - outsel1_hvt, View - schematic
// LAST TIME SAVED: Jul  3 13:08:26 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module outsel1_hvt ( out, clk, in0, in1, in2, sb, sel );
output  out;

input  clk, in0, in1, in2;

input [1:0]  sel;
input [1:0]  sb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I41 ( .A(in1), .Y(net036));
inv_hvt I40 ( .A(clk), .Y(clkb));
txgate_hvt I33 ( .in(whatever), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_hvt I_txgate1 ( .in(net036), .out(whatever), .pp(sb[0]),
     .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(whatever), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(ddr), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_hvt I38 ( .in(in2), .out(ddr), .pp(clkb), .nn(clk));
txgate_hvt I39 ( .in(in1), .out(ddr), .pp(clk), .nn(clkb));

endmodule
// Library - io, Cell - out_logic_v1, View - schematic
// LAST TIME SAVED: Jan 12 18:14:21 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module out_logic_v1 ( dout, sdo, bs_en, cbit, cbitb, ceb, clk, ddr0,
     ddr1, mode, rstio, sdi, shift, tclk, ud );
output  dout, sdo;

input  bs_en, ceb, clk, ddr0, ddr1, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbitb;
input [1:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cebdffrqn I_dff_0 ( .ceb(ceb), .clk(mux4clk), .qn(net094), .r(rstio),
     .q(sdo), .d(dd));
outsel1_hvt I_mux_func ( .clk(ddrclk), .in2(udb), .sb(cbitb[1:0]),
     .sel(cbit[1:0]), .in1(net094), .in0(dinb), .out(muxob));
nor2_hvt I_nor2 ( .A(mux4clk), .B(cbit[0]), .Y(ddrclk));
dffrckb Ireg1 ( .e(ud), .clk(mux4clk), .qn(udb), .r(rstio), .q(net44),
     .d(mux4d));
inv_hvt I171 ( .A(doutb), .Y(dout));
inv_hvt I172 ( .A(ddr0), .Y(dinb));
mux2x1_hvt I_mux_mode ( .sel(mode), .in1(udb), .in0(muxob),
     .out(doutb));
mux2x1_hvt I_mux_clk ( .in1(tclk), .in0(clk), .out(mux4clk),
     .sel(bs_en));
mux2x1_hvt I_mux_data ( .in1(sdi), .in0(ddr0), .out(dd), .sel(shift));
mux2x1_hvt I_mux_btw ( .in1(sdo), .in0(ddr1), .out(mux4d),
     .sel(bs_en));

endmodule
// Library - misc, Cell - eh_io_pup_2_new, View - schematic
// LAST TIME SAVED: Oct  6 15:01:46 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module eh_io_pup_2_new ( por_b, core_por_b, vdd_io );
output  por_b;

input  core_por_b, vdd_io;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_hvt  MP8 ( .D(net104), .B(vdd_), .G(core_por_b), .S(vdd_));
pch_hvt  M4 ( .D(por_b), .B(vdd_), .G(net92), .S(vdd_));
pch_hvt  M1 ( .D(net92), .B(vdd_), .G(net84), .S(vdd_));
pch_hvt  M0 ( .D(net84), .B(vdd_), .G(net104), .S(vdd_));
nch_hvt  M5 ( .D(por_b), .B(gnd_), .G(net92), .S(gnd_));
nch_hvt  M3 ( .D(net92), .B(gnd_), .G(net84), .S(gnd_));
nch_hvt  MN1 ( .D(net80), .B(gnd_), .G(core_por_b), .S(gnd_));
nch_hvt  M2 ( .D(net84), .B(gnd_), .G(net104), .S(gnd_));
pch_25  M6 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  MP11 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
pch_25  MP13 ( .D(net124), .B(vdd_io), .G(net145), .S(net122));
pch_25  MP12 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  M7 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  MP7 ( .D(net104), .B(vdd_), .G(net124), .S(vdd_));
pch_25  MP9 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
nch_25  MN6 ( .D(net124), .B(gnd_), .G(net145), .S(gnd_));
nch_25  MN38 ( .D(net104), .B(gnd_), .G(net124), .S(net104));
nch_25  M10 ( .D(net124), .B(gnd_), .G(net147), .S(net158));
nch_25  MN39 ( .D(net104), .B(gnd_), .G(net124), .S(net80));
nch_25  M11 ( .D(net140), .B(gnd_), .G(core_por_b), .S(gnd_));
rppolywo_m  R66 ( .MINUS(gnd_), .PLUS(net145), .BULK(gnd_));
vdd_tiehigh I96 ( .vdd_tieh(net147));
nch_na25  M15 ( .D(net154), .B(gnd_), .G(net154), .S(net150));
nch_na25  M16 ( .D(net158), .B(gnd_), .G(net158), .S(net154));
nch_na25  M17 ( .D(net162), .B(gnd_), .G(net162), .S(net166));
nch_na25  M14 ( .D(net150), .B(gnd_), .G(net150), .S(net162));
nch_na25  M18 ( .D(net166), .B(gnd_), .G(net166), .S(net140));

endmodule
// Library - io, Cell - PVSS3DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:17:04 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module PVSS3DGZ ( VSS );
input  VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - out_logic_v3, View - schematic
// LAST TIME SAVED: Jan 30 16:43:16 2008
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module out_logic_v3 ( dout, sdo, sp12, bl, bs_en, ceb, clk, ddr0, ddr1,
     mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk, ud,
     vdd_cntl, wl );
output  dout, sdo, sp12;


input  bs_en, ceb, clk, ddr0, ddr1, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;

wire  [3:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I181 ( .slfop(slfop), .cbitb(cbitb[1]), .sp12(sp12),
     .prog(prog));
cram2x2 I183 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
out_logic_v1 I_outlogic_v1 ( .ceb(ceb), .rstio(rstio), .ddr0(ddr0),
     .ddr1(ddr1), .shift(shift), .ud(ud), .clk(clk), .sdo(sdo),
     .sdi(sdi), .cbit({cbit[2], cbit[3]}), .cbitb({cbitb[2],
     cbitb[3]}), .dout(dout), .tclk(tclk), .bs_en(bs_en), .mode(mode));

endmodule
// Library - io, Cell - ioesel_hvt, View - schematic
// LAST TIME SAVED: Aug 21 18:20:13 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ioesel_hvt ( out, in0, in1, sb, sel );
output  out;

input  in0, in1;

input [1:0]  sel;
input [1:0]  sb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I38 ( .A(sel[0]), .Y(net017));
txgate_hvt I33 ( .in(mid), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_hvt I_txgate1 ( .in(in1), .out(mid), .pp(sb[0]), .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(mid), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(net017), .out(out), .pp(sel[1]), .nn(sb[1]));

endmodule
// Library - io, Cell - ioe_logic_v1, View - schematic
// LAST TIME SAVED: Jan 12 18:07:25 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ioe_logic_v1 ( outb, sdo, bs_en, cbit, cbitb, ceb, clk, din,
     mode, rstio, sdi, shift, tclk, ud );
output  outb, sdo;

input  bs_en, ceb, clk, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cebdffrqn I_dff_0 ( .ceb(ceb), .clk(net039), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_dff_1 ( .e(ud), .clk(net039), .qn(udd), .r(rstio), .q(net44),
     .d(sdo));
inv_hvt I172 ( .A(din), .Y(dinb));
mux2x1_hvt I_mux_clk ( .in1(tclk), .in0(clk), .out(net039),
     .sel(bs_en));
mux2x1_hvt I_mux_mode ( .sel(mode), .in1(udd), .in0(regmuxb),
     .out(outb));
mux2x1_hvt I_mux_data ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
ioesel_hvt I_ioe_mux2 ( .sb(cbitb[1:0]), .sel(cbit[1:0]), .in1(regb),
     .in0(dinb), .out(regmuxb));

endmodule
// Library - io, Cell - ioe_logic_v3, View - schematic
// LAST TIME SAVED: Jan 30 16:31:06 2008
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ioe_logic_v3 ( padeb, sdo, sp12, bl, bs_en, ceb, clk, din,
     hiz_b, mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk,
     ud, vdd_cntl, wl );
output  padeb, sdo, sp12;


input  bs_en, ceb, clk, din, hiz_b, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbit;

wire  [3:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[1]), .sp12(sp12),
     .prog(prog));
nand2_hvt I178 ( .A(oed), .Y(padeb), .B(hiz_b));
inv_hvt I179 ( .A(oeb), .Y(oed));
ioe_logic_v1 I_ioe_logic ( .ceb(ceb), .rstio(rstio), .cbit(cbit[3:2]),
     .cbitb(cbitb[3:2]), .outb(oeb), .bs_en(bs_en), .shift(shift),
     .ud(ud), .clk(clk), .sdo(sdo), .sdi(sdi), .din(din), .tclk(tclk),
     .mode(mode));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioe_col2rev, View - schematic
// LAST TIME SAVED: Jul 10 11:10:45 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ioe_col2rev ( dout, padeb, pado, sdo, sp12_h_l, bl, bs_en, ceb,
     hiz_b, hold, inclk, mode, outclk, padin, pgate, prog, reset,
     rstio, sdi, shift, tclk, ti, update, vdd_cntl, wl );
output  sdo;


input  bs_en, ceb, hiz_b, hold, inclk, mode, outclk, prog, rstio, sdi,
     shift, tclk, update;

output [1:0]  pado;
output [23:0]  sp12_h_l;
output [1:0]  padeb;
output [3:0]  dout;

inout [1:0]  bl;

input [1:0]  padin;
input [15:0]  vdd_cntl;
input [15:0]  reset;
input [15:0]  pgate;
input [15:0]  wl;
input [5:0]  ti;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



in_logic_v3rev I_in0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[3:2]),
     .rstio(rstio), .slfop(dout[0]), .sp12(sp12_h_l[8]), .shift(shift),
     .dout1(dout[1]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[0]), .wl(wl[3:2]), .reset(reset[3:2]),
     .sdo(s1), .sdi(s0), .pgate(pgate[3:2]), .din(padin[0]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode));
in_logic_v3rev I_in1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[13:12]),
     .rstio(rstio), .slfop(dout[3]), .sp12(sp12_h_l[14]),
     .shift(shift), .dout1(dout[3]), .ud(update), .bl(bl[1:0]),
     .prog(prog), .clk(inclk), .dout0(dout[2]), .wl(wl[13:12]),
     .reset(reset[13:12]), .sdo(s4), .sdi(s3), .pgate(pgate[13:12]),
     .din(padin[1]), .tclk(tclk), .bs_en(bs_en), .cntl(hold),
     .mode(mode));
odrv12x3 I218 ( .vdd_cntl(vdd_cntl[7:6]), .slfop({dout[1], dout[1],
     dout[1]}), .sp12({sp12_h_l[18], sp12_h_l[10], sp12_h_l[2]}),
     .bl(bl[1:0]), .wl(wl[7:6]), .reset(reset[7:6]),
     .pgate(pgate[7:6]), .prog(prog));
odrv12x3 I217 ( .vdd_cntl(vdd_cntl[9:8]), .slfop({dout[2], dout[2],
     dout[2]}), .sp12({sp12_h_l[20], sp12_h_l[12], sp12_h_l[4]}),
     .bl(bl[1:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]), .prog(prog));
out_logic_v3 I_out0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[1:0]),
     .ddr0(ti[1]), .ddr1(ti[2]), .rstio(rstio), .slfop(dout[0]),
     .sp12(sp12_h_l[0]), .dout(pado[0]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[1:0]),
     .reset(reset[1:0]), .sdo(s0), .sdi(sdi), .pgate(pgate[1:0]),
     .tclk(tclk), .bs_en(bs_en), .mode(mode));
out_logic_v3 I_out1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[11:10]),
     .ddr0(ti[4]), .ddr1(ti[5]), .rstio(rstio), .slfop(dout[3]),
     .sp12(sp12_h_l[6]), .dout(pado[1]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[11:10]),
     .reset(reset[11:10]), .sdo(s3), .sdi(s2), .pgate(pgate[11:10]),
     .tclk(tclk), .bs_en(bs_en), .mode(mode));
ioe_logic_v3 I_ioe0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[5:4]),
     .rstio(rstio), .slfop(dout[0]), .sp12(sp12_h_l[16]),
     .hiz_b(hiz_b), .padeb(padeb[0]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[5:4]),
     .reset(reset[5:4]), .sdo(s2), .sdi(s1), .pgate(pgate[5:4]),
     .din(ti[0]), .tclk(tclk), .bs_en(bs_en), .mode(mode));
ioe_logic_v3 I_ioe1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[15:14]),
     .rstio(rstio), .slfop(dout[3]), .sp12(sp12_h_l[22]),
     .hiz_b(hiz_b), .padeb(padeb[1]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[15:14]),
     .reset(reset[15:14]), .sdo(sdo), .sdi(s4), .pgate(pgate[15:14]),
     .din(ti[3]), .tclk(tclk), .bs_en(bs_en), .mode(mode));

endmodule
// Library - io, Cell - ioin_mux, View - schematic
// LAST TIME SAVED: May 18 11:01:33 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ioin_mux ( inmuxo, cbit[3], cbit[2], cbit[1], cbit[0], cbitb[3],
     cbitb[2], cbitb[1], cbitb[0], min[7:0], prog );
output  inmuxo;

input  prog;

input [0:3]  cbitb;
input [7:0]  min;
input [0:3]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I278 ( .A(net146), .Y(inmuxo));
nor2_hvt I46 ( .A(prog), .B(cbitb[3]), .Y(en));
nand2_hvt Inand2_muxo ( .A(st2), .Y(net146), .B(en));
txgate_hvt I247 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I257 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I254 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I244 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I253 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_hvt I249 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_hvt I274 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_hvt I252 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));
txgate_hvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_hvt I255 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I250 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_hvt I258 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I256 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I246 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));

endmodule
// Library - io, Cell - ioinmx1mux2rev, View - schematic
// LAST TIME SAVED: Mar  4 17:17:42 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ioinmx1mux2rev ( clk, mo, ti, bl, cdone_in, ce, ceb, in, min,
     pgate, prog, reset, spi, vdd_cntl, wl );
output  clk, ti;


input  cdone_in, ceb, prog;

output [1:0]  mo;

inout [5:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [7:0]  min;
input [1:0]  vdd_cntl;
input [1:0]  spi;
input [1:0]  reset;
input [1:0]  in;
input [11:0]  ce;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  mob;

wire  [1:0]  moo;

wire  [1:0]  r_vdd;



inv_hvt I193_1_ ( .A(moo[1]), .Y(mob[1]));
inv_hvt I193_0_ ( .A(moo[0]), .Y(mob[0]));
inv_hvt I194_1_ ( .A(mob[1]), .Y(mo[1]));
inv_hvt I194_0_ ( .A(mob[0]), .Y(mo[0]));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clk_mux12to1 I298 ( .prog(prog), .min(ce[11:0]), .clk(clk),
     .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7], cbitb[10],
     cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7], cbit[10],
     cbit[6], cbit[4]}), .cenb(ceb));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
mux2x1_hvt Iemux1_1_ ( .in1(in[1]), .in0(spi[1]), .out(moo[1]),
     .sel(cdone_in));
mux2x1_hvt Iemux1_0_ ( .in1(in[0]), .in0(spi[0]), .out(moo[0]),
     .sel(cdone_in));
ioin_mux I185 ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc, View - schematic
// LAST TIME SAVED: Aug 21 18:04:33 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  ti;
output [1:0]  spi;

inout [5:0]  bl;

input [7:0]  min2;
input [1:0]  vdd_cntl;
input [7:0]  min1;
input [1:0]  reset;
input [1:0]  padin;
input [7:0]  min0;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
nor2_hvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_hvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
inv_hvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_hvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
ioin_mux I193 ( bankcntl, {cbit[11], cbit[8], cbit[9], cbit[10]},
     {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0], prog);
ioin_mux I185 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux I186 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]}, {cbitb[5],
     cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);

endmodule
// Library - io, Cell - ioinmx2nand2inv, View - schematic
// LAST TIME SAVED: Sep 26 11:29:24 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ioinmx2nand2inv ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  ce;
input [7:0]  min0;
input [1:0]  reset;
input [7:0]  min1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
inv_hvt I181 ( .A(update), .Y(bs_enb));
nand2_hvt I180 ( .A(bs_enb), .Y(updt), .B(bs_en));
ioin_mux I185 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux I186 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]}, {cbitb[5],
     cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);

endmodule
// Library - io, Cell - sbox1mem, View - schematic
// LAST TIME SAVED: Aug 21 18:03:06 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module sbox1mem ( b, bl, l, r, t, pgate, prog, reset, vdd_cntl, wl );
inout  b, l, r, t;

input  prog;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbitb;

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox1m3to1 I232 ( .in2(r), .cb({cbitb[3], cbitb[6]}), .op(t), .in0(l),
     .in1(b), .c({cbit[3], cbit[6]}), .prog(prog));
sbox1m3to1 I230 ( .in2(r), .cb({cbitb[1], cbitb[4]}), .op(l), .in0(b),
     .in1(t), .c({cbit[1], cbit[4]}), .prog(prog));
sbox1m3to1 I226 ( .in2(r), .cb({cbitb[8], cbitb[5]}), .op(b), .in0(l),
     .in1(t), .c({cbit[8], cbit[5]}), .prog(prog));
sbox1m3to1 I231 ( .in2(b), .cb({cbitb[10], cbitb[7]}), .op(r), .in0(l),
     .in1(t), .c({cbit[10], cbit[7]}), .prog(prog));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - misc, Cell - eh_core_pup_2, View - schematic
// LAST TIME SAVED: Jul 11 11:51:16 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module eh_core_pup_2 ( por_b );
output  por_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo  R10 ( .MINUS(net130), .PLUS(net109));
rppolywo  R12 ( .MINUS(net154), .PLUS(net157));
rppolywo  R6 ( .MINUS(out_1), .PLUS(net124));
rppolywo  R9 ( .MINUS(net118), .PLUS(net130));
rppolywo  R15 ( .MINUS(net166), .PLUS(div_1));
rppolywo  R13 ( .MINUS(net157), .PLUS(net145));
rppolywo  R1 ( .MINUS(net068), .PLUS(net048));
rppolywo  R2 ( .MINUS(net067), .PLUS(net068));
rppolywo  R4 ( .MINUS(net142), .PLUS(net148));
rppolywo  R5 ( .MINUS(div_1), .PLUS(net142));
rppolywo  R41 ( .MINUS(net039), .PLUS(net042));
rppolywo  R40 ( .MINUS(net042), .PLUS(vdd_));
rppolywo  R11 ( .MINUS(net109), .PLUS(net154));
rppolywo  R0 ( .MINUS(net048), .PLUS(net039));
rppolywo  R8 ( .MINUS(net127), .PLUS(net118));
rppolywo  R14 ( .MINUS(net145), .PLUS(net166));
rppolywo  R3 ( .MINUS(net148), .PLUS(net067));
rppolywo  R7 ( .MINUS(net124), .PLUS(net127));
nch_hvt  M0 ( .D(out_1), .B(gnd_), .G(div_1), .S(gnd_));
nch_hvt  M2 ( .D(out_1), .B(gnd_), .G(out_2), .S(gnd_));
nch_hvt  M6 ( .D(gnd_), .B(gnd_), .G(out_2), .S(gnd_));
inv_hvt I11 ( .A(out_4), .Y(net193));
inv_hvt I2 ( .A(out_3), .Y(out_4));
inv_hvt I7 ( .A(out_1), .Y(out_2));
inv_hvt I9 ( .A(out_2), .Y(out_3));
inv_hvt I6 ( .A(net193), .Y(por_b));

endmodule
// Library - io, Cell - sbox1_colbdlc_rev, View - schematic
// LAST TIME SAVED: Jul 10 10:35:15 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module sbox1_colbdlc_rev ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  pado;
output [1:0]  spi_ss_in_b;
output [5:0]  ti;
output [1:0]  padeb;

inout [5:0]  bl;
inout [3:0]  l;
inout [3:0]  sp4_v_b;
inout [3:0]  r;
inout [3:0]  t_mid;

input [1:0]  padin;
input [7:0]  ceb_in;
input [1:0]  spiout;
input [11:0]  clk_in;
input [7:0]  min0;
input [1:0]  oeb;
input [7:0]  min1;
input [1:0]  out;
input [7:0]  min3;
input [7:0]  min6;
input [1:0]  spioeb;
input [7:0]  min4;
input [7:0]  min5;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [11:0]  inclk_in;
input [7:0]  min2;
input [15:0]  reset;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ioinmx1mux2rev I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .in(out[1:0]), .ti(ti[2]), .min(min2[7:0]), .spi(spiout[1:0]),
     .wl(wl[9:8]), .reset(reset[9:8]), .pgate(pgate[9:8]),
     .cdone_in(cdone_in), .mo(pado[1:0]));
ioinmx1mux2rev I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .in(oeb[1:0]), .ti(ti[5]), .min(min5[7:0]), .spi(spioeb[1:0]),
     .wl(wl[15:14]), .reset(reset[15:14]), .pgate(pgate[15:14]),
     .cdone_in(cdone_in), .mo(padeb[1:0]));
ioinmx2nor2invx2bdlc I5 ( .vdd_cntl(vdd_cntl[5:4]), .min2(min6[7:0]),
     .bankcntl(fabric_out), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx2nand2inv I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - io, Cell - io_odrv4x5, View - schematic
// LAST TIME SAVED: Aug 21 17:59:07 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module io_odrv4x5 ( cbit, sp4_out, bl, pgate, prog,
     reset, slfop, vdd_cntl, wl );


input  prog, slfop;

output [4:0]  sp4_out;
output [7:5]  cbit;

inout [3:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
supply0 gnd_;
supply1 vdd_;

// Buses in the design

wire  [7:0]  cbitb;

wire  [1:0]  r_vdd;

wire [7:0] cbit_int;
assign cbit[7:5] = cbit_int[7:5];


pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv4 I_odrv_4_ ( .cbitb(cbitb[4]), .sp4(sp4_out[4]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_3_ ( .cbitb(cbitb[3]), .sp4(sp4_out[3]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_2_ ( .cbitb(cbitb[2]), .sp4(sp4_out[2]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_1_ ( .cbitb(cbitb[1]), .sp4(sp4_out[1]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_0_ ( .cbitb(cbitb[0]), .sp4(sp4_out[0]), .slfop(slfop),
     .prog(prog));
cram2x2 Icram2x2_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset[1:0]), .q(cbit_int[7:4]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));
cram2x2 Icram2x2_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset[1:0]), .q(cbit_int[3:0]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - io_col_odrv4_x40bare, View - schematic
// LAST TIME SAVED: Jul 31 17:45:40 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module io_col_odrv4_x40bare ( cf, bl, sp4_h_l,
     sp4_v_b, dout0, dout1,
     pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [23:0]  cf;

inout [3:0]  bl;
inout [15:0]  sp4_v_b;
inout [47:0]  sp4_h_l;

input [0:1]  dout0;
input [0:1]  dout1;
input [15:0]  pgate;
input [15:0]  wl;
input [15:0]  reset;
input [15:0]  vdd_cntl;
supply0 gnd_;
supply1 vdd_;



io_odrv4x5 I218 ( cf[20:18], {sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6]}, bl[3:0], pgate[13:12], prog,
     reset[13:12], dout1[1], vdd_cntl[13:12], wl[13:12]);
io_odrv4x5 I217 ( cf[14:12], {sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4]}, bl[3:0], pgate[9:8], prog, reset[9:8],
     dout0[1], vdd_cntl[9:8], wl[9:8]);
io_odrv4x5 I_odrv_4x5_7 ( cf[23:21], {sp4_v_b[15], sp4_v_b[11],
     sp4_v_b[7], sp4_v_b[3], sp4_h_l[46]}, bl[3:0], pgate[15:14], prog,
     reset[15:14], dout1[1], vdd_cntl[15:14], wl[15:14]);
io_odrv4x5 I220 ( cf[11:9], {sp4_v_b[13], sp4_v_b[9], sp4_v_b[5],
     sp4_v_b[1], sp4_h_l[42]}, bl[3:0], pgate[7:6], prog, reset[7:6],
     dout1[0], vdd_cntl[7:6], wl[7:6]);
io_odrv4x5 I221 ( cf[8:6], {sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2]}, bl[3:0], pgate[5:4], prog, reset[5:4],
     dout1[0], vdd_cntl[5:4], wl[5:4]);
io_odrv4x5 I_odrv_4x5_0 ( cf[2:0], {sp4_h_l[32], sp4_h_l[24],
     sp4_h_l[16], sp4_h_l[8], sp4_h_l[0]}, bl[3:0], pgate[1:0], prog,
     reset[1:0], dout0[0], vdd_cntl[1:0], wl[1:0]);
io_odrv4x5 I223 ( cf[5:3], {sp4_v_b[12], sp4_v_b[8], sp4_v_b[4],
     sp4_v_b[0], sp4_h_l[40]}, bl[3:0], pgate[3:2], prog, reset[3:2],
     dout0[0], vdd_cntl[3:2], wl[3:2]);
io_odrv4x5 I215 ( cf[17:15], {sp4_v_b[14], sp4_v_b[10], sp4_v_b[6],
     sp4_v_b[2], sp4_h_l[44]}, bl[3:0], pgate[11:10], prog,
     reset[11:10], dout0[1], vdd_cntl[11:10], wl[11:10]);

endmodule
// Library - io, Cell - io_gmux_x2, View - schematic
// LAST TIME SAVED: Jan  7 13:58:08 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module io_gmux_x2 ( .cbit_colcntl({cbit[11], cbit[9]}), gout, bl, min0,
     min1, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [1:0]  gout;
output [11:0]  cbit;

inout [5:0]  bl;

input [1:0]  reset;
input [15:0]  min1;
input [1:0]  wl;
input [15:0]  min0;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux Ig_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux Ig_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - io, Cell - io_gmux_x16bare, View - schematic
// LAST TIME SAVED: Feb 19 09:24:32 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module io_gmux_x16bare ( cbit_colcntl, lc_trk_g0, lc_trk_g1, bl, min0,
     min1, min2, min3, min4, min5, min6, min7, min8, min9, min10,
     min11, min12, min13, min14, min15, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [7:0]  cbit_colcntl;
output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;

inout [5:0]  bl;

input [15:0]  min0;
input [15:0]  min9;
input [15:0]  min13;
input [15:0]  min10;
input [15:0]  min7;
input [15:0]  min1;
input [15:0]  min12;
input [15:0]  min2;
input [15:0]  min3;
input [15:0]  min11;
input [15:0]  min8;
input [15:0]  min5;
input [15:0]  min4;
input [15:0]  reset;
input [15:0]  min15;
input [15:0]  pgate;
input [15:0]  min6;
input [15:0]  wl;
input [15:0]  vdd_cntl;
input [15:0]  min14;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net132;

wire  [0:1]  net122;

wire  [0:1]  net182;

wire  [0:1]  net112;



io_gmux_x2 Iio_gmux4 ( .cbit_colcntl(net112[0:1]),
     .vdd_cntl(vdd_cntl[9:8]), .bl(bl[5:0]), .min0(min8[15:0]),
     .gout(lc_trk_g1[1:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]), .min1(min9[15:0]), .prog(prog));
io_gmux_x2 Iio_gmux5 ( .cbit_colcntl(net122[0:1]),
     .vdd_cntl(vdd_cntl[11:10]), .bl(bl[5:0]), .min0(min10[15:0]),
     .gout(lc_trk_g1[3:2]), .wl(wl[11:10]), .reset(reset[11:10]),
     .pgate(pgate[11:10]), .min1(min11[15:0]), .prog(prog));
io_gmux_x2 Iio_gmux6 ( .cbit_colcntl(net132[0:1]),
     .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .min0(min12[15:0]),
     .gout(lc_trk_g1[5:4]), .wl(wl[13:12]), .reset(reset[13:12]),
     .pgate(pgate[13:12]), .min1(min13[15:0]), .prog(prog));
io_gmux_x2 Iio_gmux1 ( .cbit_colcntl(cbit_colcntl[3:2]),
     .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .min0(min2[15:0]),
     .gout(lc_trk_g0[3:2]), .wl(wl[3:2]), .reset(reset[3:2]),
     .pgate(pgate[3:2]), .min1(min3[15:0]), .prog(prog));
io_gmux_x2 Iio_gmux0 ( .cbit_colcntl(cbit_colcntl[1:0]),
     .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .min0(min0[15:0]),
     .gout(lc_trk_g0[1:0]), .wl(wl[1:0]), .reset(reset[1:0]),
     .pgate(pgate[1:0]), .min1(min1[15:0]), .prog(prog));
io_gmux_x2 Iio_gmux2 ( .cbit_colcntl(cbit_colcntl[5:4]),
     .vdd_cntl(vdd_cntl[5:4]), .bl(bl[5:0]), .min0(min4[15:0]),
     .gout(lc_trk_g0[5:4]), .wl(wl[5:4]), .reset(reset[5:4]),
     .pgate(pgate[5:4]), .min1(min5[15:0]), .prog(prog));
io_gmux_x2 Iio_gmux3 ( .cbit_colcntl(cbit_colcntl[7:6]),
     .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .min0(min6[15:0]),
     .gout(lc_trk_g0[7:6]), .wl(wl[7:6]), .reset(reset[7:6]),
     .pgate(pgate[7:6]), .min1(min7[15:0]), .prog(prog));
io_gmux_x2 Iio_gmux7 ( .cbit_colcntl(net182[0:1]),
     .vdd_cntl(vdd_cntl[15:14]), .bl(bl[5:0]), .min0(min14[15:0]),
     .gout(lc_trk_g1[7:6]), .wl(wl[15:14]), .reset(reset[15:14]),
     .pgate(pgate[15:14]), .min1(min15[15:0]), .prog(prog));

endmodule
// Library - io, Cell - io_col4_LFT_rev, View - schematic
// LAST TIME SAVED: Apr 28 16:05:00 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module io_col4_LFT_rev ( cbit_colcntl, cf, fabric_out, padeb, pado,
     sdo, slf_op, spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l,
     bnl_op, bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op,
     mode, padin, pgate, prog, r, reset, sdi, shift, spioeb, spiout,
     tclk, tnl_op, update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [7:0]  cbit_colcntl;
output [1:0]  padeb;
output [23:0]  cf;
output [3:0]  slf_op;
output [1:0]  spi_ss_in_b;
output [1:0]  pado;

inout [15:0]  sp4_v_t;
inout [17:0]  bl;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;

input [1:0]  spiout;
input [15:0]  wl;
input [15:0]  vdd_cntl;
input [15:0]  reset;
input [15:0]  pgate;
input [1:0]  spioeb;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  glb_netwk;
input [1:0]  padin;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



ioe_col2rev I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .dout(slf_op[3:0]), .outclk(outclk), .hold(hold),
     .rstio(r), .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]}), .reset({reset[14], reset[15], reset[12], reset[13],
     reset[10], reset[11], reset[8], reset[9], reset[6], reset[7],
     reset[4], reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net127), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));
sbox1_colbdlc_rev Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net127));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net127));
rm7  R14_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7  R14_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7  R14_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7  R14_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7  R14_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7  R14_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7  R14_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7  R14_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7  R14_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7  R14_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7  R14_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7  R14_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7  R14_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7  R14_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7  R14_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7  R14_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net127, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .cbit_colcntl(cbit_colcntl[7:0]),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min7({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}), .min5({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14], wl[15],
     wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4],
     wl[5], wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .prog(net127),
     .lc_trk_g1(lc_trk_g1[7:0]));

endmodule
// Library - leafcell, Cell - clk_colbuf1k, View - schematic
// LAST TIME SAVED: Feb 12 17:34:53 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module clk_colbuf1k ( clko, cbit, clki );
output  clko;

input  cbit, clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(clko), .B(gnd_), .G(clkb), .S(net7));
nch_hvt  M2 ( .D(net7), .B(gnd_), .G(cbit), .S(gnd_));
pch_hvt  M0 ( .D(clko), .B(vdd_), .G(clkb), .S(vdd_));
nand2_hvt I_nand2_hvt ( .A(clki), .Y(clkb), .B(cbit));

endmodule
// Library - leafcell, Cell - clk_colbuf1kx8, View - schematic
// LAST TIME SAVED: Apr 27 11:45:11 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module clk_colbuf1kx8 ( col_clk, clk_in, colbuf_cntl );


output [7:0]  col_clk;

input [7:0]  clk_in;
input [7:0]  colbuf_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clk_colbuf1k I_colbuf1k_7_ ( .clki(clk_in[7]), .clko(col_clk[7]),
     .cbit(colbuf_cntl[7]));
clk_colbuf1k I_colbuf1k_6_ ( .clki(clk_in[6]), .clko(col_clk[6]),
     .cbit(colbuf_cntl[6]));
clk_colbuf1k I_colbuf1k_5_ ( .clki(clk_in[5]), .clko(col_clk[5]),
     .cbit(colbuf_cntl[5]));
clk_colbuf1k I_colbuf1k_4_ ( .clki(clk_in[4]), .clko(col_clk[4]),
     .cbit(colbuf_cntl[4]));
clk_colbuf1k I_colbuf1k_3_ ( .clki(clk_in[3]), .clko(col_clk[3]),
     .cbit(colbuf_cntl[3]));
clk_colbuf1k I_colbuf1k_2_ ( .clki(clk_in[2]), .clko(col_clk[2]),
     .cbit(colbuf_cntl[2]));
clk_colbuf1k I_colbuf1k_1_ ( .clki(clk_in[1]), .clko(col_clk[1]),
     .cbit(colbuf_cntl[1]));
clk_colbuf1k I_colbuf1k_0_ ( .clki(clk_in[0]), .clko(col_clk[0]),
     .cbit(colbuf_cntl[0]));

endmodule
// Library - leafcell, Cell - ice1f_array_LFT_IO_bot14io, View -
//schematic
// LAST TIME SAVED: Aug 14 12:00:37 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ice1f_array_LFT_IO_bot14io ( cf_l, fabric_out_01, fabric_out_02,
     fabric_out_03, fabric_out_04, fabric_out_05, fabric_out_06,
     fabric_out_07, fabric_out_08, padeb, pado, sdo, slf_op_00_01,
     slf_op_00_02, slf_op_00_03, slf_op_00_04, slf_op_00_05,
     slf_op_00_06, slf_op_00_07, slf_op_00_08, spi_ss_in_b,
     SP4_h_l_00_01, SP4_h_l_00_02, SP4_h_l_00_03, SP4_h_l_00_04,
     SP4_h_l_00_05, SP4_h_l_00_06, SP4_h_l_00_07, SP4_h_l_00_08,
     SP12_h_l_00_01, SP12_h_l_00_02, SP12_h_l_00_03, SP12_h_l_00_04,
     SP12_h_l_00_05, SP12_h_l_00_06, SP12_h_l_00_07, SP12_h_l_00_08,
     bl, pgate, reset_b, sp4_v_b_00_01, sp4_v_t_00_08, vdd_cntl, wl,
     bnl_op_00_01, bs_en, cdone_in, ceb, glb_netwk_col, hiz_b, hold,
     mode, padin, prog, r, rgt_op_00_01, rgt_op_00_02, rgt_op_00_03,
     rgt_op_00_04, rgt_op_00_05, rgt_op_00_06, rgt_op_00_07,
     rgt_op_00_08, sdi, shift, spioeb, spiout, tclk, tnl_op_00_08,
     update );
output  fabric_out_01, fabric_out_02, fabric_out_03, fabric_out_04,
     fabric_out_05, fabric_out_06, fabric_out_07, fabric_out_08, sdo;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_00_07;
output [3:0]  slf_op_00_04;
output [3:0]  slf_op_00_03;
output [3:0]  slf_op_00_06;
output [3:0]  slf_op_00_01;
output [3:0]  slf_op_00_08;
output [3:0]  slf_op_00_02;
output [3:0]  slf_op_00_05;
output [13:0]  padeb;
output [191:0]  cf_l;
output [15:0]  spi_ss_in_b;
output [13:0]  pado;

inout [23:0]  SP12_h_l_00_03;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_00_06;
inout [15:0]  sp4_v_b_00_01;
inout [23:0]  SP12_h_l_00_06;
inout [23:0]  SP12_h_l_00_08;
inout [47:0]  SP4_h_l_00_02;
inout [23:0]  SP12_h_l_00_01;
inout [23:0]  SP12_h_l_00_04;
inout [47:0]  SP4_h_l_00_05;
inout [47:0]  SP4_h_l_00_08;
inout [15:0]  sp4_v_t_00_08;
inout [23:0]  SP12_h_l_00_07;
inout [47:0]  SP4_h_l_00_07;
inout [23:0]  SP12_h_l_00_05;
inout [47:0]  SP4_h_l_00_01;
inout [23:0]  SP12_h_l_00_02;
inout [47:0]  SP4_h_l_00_04;
inout [47:0]  SP4_h_l_00_03;
inout [127:0]  reset_b;
inout [127:0]  vdd_cntl;
inout [127:0]  pgate;
inout [127:0]  wl;

input [7:0]  rgt_op_00_07;
input [7:0]  rgt_op_00_02;
input [7:0]  glb_netwk_col;
input [7:0]  bnl_op_00_01;
input [7:0]  rgt_op_00_05;
input [7:0]  rgt_op_00_03;
input [7:0]  rgt_op_00_08;
input [7:0]  tnl_op_00_08;
input [7:0]  rgt_op_00_04;
input [7:0]  rgt_op_00_06;
input [7:0]  rgt_op_00_01;
input [15:0]  spiout;
input [13:0]  padin;
input [15:0]  spioeb;
input [8:1]  cdone_in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net601;

wire  [7:0]  glb_netwk_b;

wire  [7:0]  colbuf_cntl_b;

wire  [7:0]  colbuf_cntl_t;

wire  [7:0]  glb_netwk_t;

wire  [0:1]  net383;

wire  [0:7]  net634;

wire  [0:15]  net385;

wire  [0:15]  net421;

wire  [0:1]  net628;

wire  [0:15]  net457;

wire  [0:15]  net493;

wire  [0:7]  net631;

wire  [0:15]  net529;

wire  [0:7]  net633;

wire  [15:0]  colbuf_cntl;

wire  [0:15]  net565;

wire  [0:7]  net636;



io_col4_LFT_rev I_io_00_08 ( .cbit_colcntl(net634[0:7]), .ceb(ceb),
     .sdo(net371), .sdi(sdi), .spiout(spiout[15:14]),
     .cdone_in(cdone_in[8]), .spioeb(spioeb[15:14]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[13:12]), .pado(pado[13:12]),
     .padeb(padeb[13:12]), .sp4_v_t(sp4_v_t_00_08[15:0]),
     .sp4_h_l(SP4_h_l_00_08[47:0]), .sp12_h_l(SP12_h_l_00_08[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[15:14]),
     .tnl_op(tnl_op_00_08[7:0]), .lft_op(rgt_op_00_08[7:0]),
     .bnl_op(rgt_op_00_07[7:0]), .pgate(pgate[127:112]),
     .reset(reset_b[127:112]), .sp4_v_b(net385[0:15]),
     .wl(wl[127:112]), .cf(cf_l[191:168]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[127:112]), .slf_op(slf_op_00_08[3:0]),
     .glb_netwk(glb_netwk_t[7:0]), .hold(hold),
     .fabric_out(fabric_out_08));
io_col4_LFT_rev I_io_00_07 ( .cbit_colcntl(net631[0:7]), .ceb(ceb),
     .sdo(net443), .sdi(net371), .spiout(spiout[13:12]),
     .cdone_in(cdone_in[7]), .spioeb(spioeb[13:12]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(net383[0:1]), .pado(net383[0:1]),
     .padeb(net628[0:1]), .sp4_v_t(net385[0:15]),
     .sp4_h_l(SP4_h_l_00_07[47:0]), .sp12_h_l(SP12_h_l_00_07[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[13:12]),
     .tnl_op(rgt_op_00_08[7:0]), .lft_op(rgt_op_00_07[7:0]),
     .bnl_op(rgt_op_00_06[7:0]), .pgate(pgate[111:96]),
     .reset(reset_b[111:96]), .sp4_v_b(net457[0:15]), .wl(wl[111:96]),
     .cf(cf_l[167:144]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_00_07[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_07));
io_col4_LFT_rev I_io_00_05 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net587), .sdi(net407), .spiout(spiout[9:8]),
     .cdone_in(cdone_in[5]), .spioeb(spioeb[9:8]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[9:8]), .pado(pado[9:8]),
     .padeb(padeb[9:8]), .sp4_v_t(net421[0:15]),
     .sp4_h_l(SP4_h_l_00_05[47:0]), .sp12_h_l(SP12_h_l_00_05[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[9:8]),
     .tnl_op(rgt_op_00_06[7:0]), .lft_op(rgt_op_00_05[7:0]),
     .bnl_op(rgt_op_00_04[7:0]), .pgate(pgate[79:64]),
     .reset(reset_b[79:64]), .sp4_v_b(net601[0:15]), .wl(wl[79:64]),
     .cf(cf_l[119:96]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_00_05[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_05));
io_col4_LFT_rev I_io_00_06 ( .cbit_colcntl(net633[0:7]), .ceb(ceb),
     .sdo(net407), .sdi(net443), .spiout(spiout[11:10]),
     .cdone_in(cdone_in[6]), .spioeb(spioeb[11:10]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[11:10]), .pado(pado[11:10]),
     .padeb(padeb[11:10]), .sp4_v_t(net457[0:15]),
     .sp4_h_l(SP4_h_l_00_06[47:0]), .sp12_h_l(SP12_h_l_00_06[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[11:10]),
     .tnl_op(rgt_op_00_07[7:0]), .lft_op(rgt_op_00_06[7:0]),
     .bnl_op(rgt_op_00_05[7:0]), .pgate(pgate[95:80]),
     .reset(reset_b[95:80]), .sp4_v_b(net421[0:15]), .wl(wl[95:80]),
     .cf(cf_l[143:120]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_00_06[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_06));
io_col4_LFT_rev I_io_00_02 ( .cbit_colcntl(colbuf_cntl[15:8]),
     .ceb(ceb), .sdo(net515), .sdi(net479), .spiout(spiout[3:2]),
     .cdone_in(cdone_in[2]), .spioeb(spioeb[3:2]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[3:2]), .pado(pado[3:2]),
     .padeb(padeb[3:2]), .sp4_v_t(net493[0:15]),
     .sp4_h_l(SP4_h_l_00_02[47:0]), .sp12_h_l(SP12_h_l_00_02[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[3:2]),
     .tnl_op(rgt_op_00_03[7:0]), .lft_op(rgt_op_00_02[7:0]),
     .bnl_op(rgt_op_00_01[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b(net529[0:15]), .wl(wl[31:16]),
     .cf(cf_l[47:24]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_00_02[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_02));
io_col4_LFT_rev I_io_00_01 ( .cbit_colcntl(colbuf_cntl[7:0]),
     .ceb(ceb), .sdo(sdo), .sdi(net515), .spiout(spiout[1:0]),
     .cdone_in(cdone_in[1]), .spioeb(spioeb[1:0]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .sp4_v_t(net529[0:15]),
     .sp4_h_l(SP4_h_l_00_01[47:0]), .sp12_h_l(SP12_h_l_00_01[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[1:0]),
     .tnl_op(rgt_op_00_02[7:0]), .lft_op(rgt_op_00_01[7:0]),
     .bnl_op(bnl_op_00_01[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(sp4_v_b_00_01[15:0]),
     .wl(wl[15:0]), .cf(cf_l[23:0]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_00_01[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold),
     .fabric_out(fabric_out_01));
io_col4_LFT_rev I_io_00_03 ( .cbit_colcntl(net636[0:7]), .ceb(ceb),
     .sdo(net479), .sdi(net551), .spiout(spiout[5:4]),
     .cdone_in(cdone_in[3]), .spioeb(spioeb[5:4]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[5:4]), .pado(pado[5:4]),
     .padeb(padeb[5:4]), .sp4_v_t(net565[0:15]),
     .sp4_h_l(SP4_h_l_00_03[47:0]), .sp12_h_l(SP12_h_l_00_03[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[5:4]),
     .tnl_op(rgt_op_00_04[7:0]), .lft_op(rgt_op_00_03[7:0]),
     .bnl_op(rgt_op_00_02[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b(net493[0:15]), .wl(wl[47:32]),
     .cf(cf_l[71:48]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_00_03[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_03));
io_col4_LFT_rev I_io_00_04 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net551), .sdi(net587), .spiout(spiout[7:6]),
     .cdone_in(cdone_in[4]), .spioeb(spioeb[7:6]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[7:6]), .pado(pado[7:6]),
     .padeb(padeb[7:6]), .sp4_v_t(net601[0:15]),
     .sp4_h_l(SP4_h_l_00_04[47:0]), .sp12_h_l(SP12_h_l_00_04[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[7:6]),
     .tnl_op(rgt_op_00_05[7:0]), .lft_op(rgt_op_00_04[7:0]),
     .bnl_op(rgt_op_00_03[7:0]), .pgate(pgate[63:48]),
     .reset(reset_b[63:48]), .sp4_v_b(net565[0:15]), .wl(wl[63:48]),
     .cf(cf_l[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_00_04[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_04));
clk_colbuf1kx8 I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_colbuf1kx8 I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - io, Cell - io_col4_BOT_rev, View - schematic
// LAST TIME SAVED: Apr 28 16:01:05 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module io_col4_BOT_rev ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  padeb;
output [1:0]  pado;
output [23:0]  cf;
output [3:0]  slf_op;
output [1:0]  spi_ss_in_b;

inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;
inout [17:0]  bl;
inout [47:0]  sp4_h_l;
inout [23:0]  sp12_h_l;

input [1:0]  padin;
input [1:0]  spioeb;
input [1:0]  spiout;
input [15:0]  reset;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  glb_netwk;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net0140;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [1:0]  oenm;

wire  [5:0]  ti;

wire  [3:0]  t_mid;

wire  [1:0]  om;



ioe_col2rev I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .dout(slf_op[3:0]), .outclk(outclk), .hold(hold),
     .rstio(r), .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]}), .reset({reset[14], reset[15], reset[12], reset[13],
     reset[10], reset[11], reset[8], reset[9], reset[6], reset[7],
     reset[4], reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net0214), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));
sbox1_colbdlc_rev Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net0214));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net0214));
rm6  R14_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6  R14_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6  R14_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6  R14_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6  R14_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6  R14_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6  R14_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6  R14_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6  R14_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6  R14_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6  R14_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6  R14_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6  R14_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6  R14_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6  R14_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6  R14_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net0214, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .cbit_colcntl(net0140[0:7]),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min7({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}), .min5({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14], wl[15],
     wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4],
     wl[5], wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .prog(net0214),
     .lc_trk_g1(lc_trk_g1[7:0]));

endmodule
// Library - misc, Cell - SMC_CORE_POR_right, View - schematic
// LAST TIME SAVED: Aug 14 14:25:50 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module SMC_CORE_POR_right ( core_por_b, smc_por_b, creset_b,
     smc_core_por_bottom1, smc_core_por_bottom2, vddio_rightbank );
output  core_por_b, smc_por_b;

input  creset_b, smc_core_por_bottom1, smc_core_por_bottom2,
     vddio_rightbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I6 ( .A(net026), .Y(net021), .B(creset_b));
eh_io_pup_2_new I0 ( .vdd_io(vddio_rightbank), .core_por_b(net026),
     .por_b(net3));
eh_core_pup_2 I1 ( .por_b(net026));
nand4_hvt I2 ( .D(core_por_b), .C(smc_core_por_bottom2), .A(net3),
     .Y(net04), .B(smc_core_por_bottom1));
inv_hvt I7 ( .A(net021), .Y(core_por_b));
inv_hvt I3 ( .A(net04), .Y(smc_por_b));

endmodule
// Library - leafcell, Cell - tckbufx16, View - schematic
// LAST TIME SAVED: Jan 31 14:34:05 2008
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module tckbufx16 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - bram_bufferx4x6, View - schematic
// LAST TIME SAVED: Sep 15 13:53:57 2008
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module bram_bufferx4x6 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I4 ( .in(d1), .out(d2));
bram_bufferx4 I5 ( .in(d2), .out(d3));
bram_bufferx4 I6 ( .in(d3), .out(d4));
bram_bufferx4 I7 ( .in(d4), .out(out));
bram_bufferx4 I3 ( .in(d0), .out(d1));
bram_bufferx4 I0 ( .in(in), .out(d0));

endmodule
// Library - leafcell, Cell - lowla_modified, View - schematic
// LAST TIME SAVED: Sep 15 13:19:27 2008
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module lowla_modified ( lao, clk, min );
output  lao;

input  clk, min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I289 ( .A(net29), .Y(lao));
inv_hvt I290 ( .A(st2), .Y(net29));
inv_hvt I_inv ( .A(clk), .Y(cbitb));
inv_hvt I_inv3 ( .A(cbitb), .Y(clkd));
txgate_hvt I249 ( .in(lao), .out(st2), .pp(cbitb), .nn(clkd));
txgate_hvt I248 ( .in(min), .out(st2), .pp(clkd), .nn(cbitb));

endmodule
// Library - leafcell, Cell - scanbuf1f, View - schematic
// LAST TIME SAVED: Jun 10 18:32:28 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module scanbuf1f ( bs_en_o, ceb_o, hiz_b_o, mode_o, r_o, sdo, shift_o,
     tclk_o, update_o, bs_en_i, ceb_i, hiz_b_i, mode_i, r_i, sdi,
     shift_i, tclk_i, update_i );
output  bs_en_o, ceb_o, hiz_b_o, mode_o, r_o, sdo, shift_o, tclk_o,
     update_o;

input  bs_en_i, ceb_i, hiz_b_i, mode_i, r_i, sdi, shift_i, tclk_i,
     update_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



tckbufx16 I_tclkbuf ( .in(tclk_i), .out(tclk_o));
bram_bufferx4 I_bs_enbuf ( .in(bs_en_i), .out(bs_en_o));
bram_bufferx4 I_cebbuf ( .in(ceb_i), .out(ceb_o));
bram_bufferx4 I_modebuf ( .in(mode_i), .out(mode_o));
bram_bufferx4 I_hiz_bbuf ( .in(hiz_b_i), .out(hiz_b_o));
bram_bufferx4 I_updatebuf ( .in(update_i), .out(update_o));
bram_bufferx4 I_shiftbuf ( .in(shift_i), .out(shift_o));
bram_bufferx4 I_rbuf ( .in(r_i), .out(r_o));
bram_bufferx4x6 I_sdibuf ( .in(sdi), .out(sdi_2));
lowla_modified I_lowla ( .clk(tclk_i), .min(sdi_2), .lao(sdo));

endmodule
// Library - leafcell, Cell - ice1f_array_BOT_IO_lft12io, View -
//schematic
// LAST TIME SAVED: Jul 22 08:44:03 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module ice1f_array_BOT_IO_lft12io ( bs_en_o, ceb_o, cf_bot_l,
     fabric_out_05_00, fabric_out_06_00, hiz_b_o, mode_o, padeb_b_l,
     pado_b_l, r_o, sdo, shift_o, slf_op_01_00, slf_op_02_00,
     slf_op_03_00, slf_op_04_00, slf_op_05_00, slf_op_06_00, tclk_o,
     update_o, bl_01, bl_02, bl_03, bl_04, bl_05, bl_06, sp4_h_l_01_00,
     sp4_h_r_06_00, sp4_v_b_01_00, sp4_v_b_02_00, sp4_v_b_03_00,
     sp4_v_b_04_00, sp4_v_b_05_00, sp4_v_b_06_00, sp12_v_b_01_00,
     sp12_v_b_02_00, sp12_v_b_03_00, sp12_v_b_04_00, sp12_v_b_05_00,
     sp12_v_b_06_00, bnl_op_01_00, bs_en_i, ceb_i, glb_net_01,
     glb_net_02, glb_net_03, glb_net_04, glb_net_05, glb_net_06,
     hiz_b_i, hold_b_l, lft_op_01_00, lft_op_02_00, lft_op_03_00,
     lft_op_04_00, lft_op_05_00, lft_op_06_00, mode_i, padin_b_l,
     pgate_l, prog, r_i, reset_l, sdi, shift_i, tclk_i, tiegnd, tievdd,
     tnr_op_06_00, update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_05_00, fabric_out_06_00, hiz_b_o,
     mode_o, r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_b_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, tiegnd, tievdd, update_i;

output [3:0]  slf_op_04_00;
output [3:0]  slf_op_03_00;
output [3:0]  slf_op_01_00;
output [3:0]  slf_op_05_00;
output [3:0]  slf_op_06_00;
output [11:0]  padeb_b_l;
output [11:0]  pado_b_l;
output [143:0]  cf_bot_l;
output [3:0]  slf_op_02_00;

inout [47:0]  sp4_v_b_03_00;
inout [47:0]  sp4_v_b_06_00;
inout [23:0]  sp12_v_b_06_00;
inout [23:0]  sp12_v_b_04_00;
inout [23:0]  sp12_v_b_02_00;
inout [15:0]  sp4_h_r_06_00;
inout [47:0]  sp4_v_b_04_00;
inout [23:0]  sp12_v_b_01_00;
inout [47:0]  sp4_v_b_01_00;
inout [47:0]  sp4_v_b_02_00;
inout [23:0]  sp12_v_b_05_00;
inout [41:0]  bl_03;
inout [53:0]  bl_06;
inout [53:0]  bl_04;
inout [53:0]  bl_05;
inout [53:0]  bl_02;
inout [47:0]  sp4_v_b_05_00;
inout [15:0]  sp4_h_l_01_00;
inout [23:0]  sp12_v_b_03_00;
inout [53:0]  bl_01;

input [15:0]  wl_l;
input [7:0]  glb_net_04;
input [7:0]  lft_op_06_00;
input [7:0]  bnl_op_01_00;
input [15:0]  pgate_l;
input [7:0]  lft_op_02_00;
input [7:0]  tnr_op_06_00;
input [7:0]  lft_op_03_00;
input [7:0]  glb_net_05;
input [7:0]  glb_net_01;
input [7:0]  glb_net_03;
input [15:0]  vdd_cntl_l;
input [7:0]  lft_op_05_00;
input [11:0]  padin_b_l;
input [7:0]  glb_net_06;
input [7:0]  lft_op_04_00;
input [7:0]  glb_net_02;
input [15:0]  reset_l;
input [7:0]  lft_op_01_00;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net364;

wire  [0:15]  net329;

wire  [0:1]  net497;

wire  [0:1]  net492;

wire  [0:15]  net399;

wire  [0:1]  net502;

wire  [0:1]  net501;

wire  [0:15]  net434;

wire  [0:1]  net473;

wire  [0:1]  net333;

wire  [0:15]  net294;



io_col4_BOT_rev I_io_t01 ( .sdo(net278), .sdi(sdi), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .sp4_v_t(sp4_h_l_01_00[15:0]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_b_l[1:0]), .pado(pado_b_l[1:0]),
     .padeb(padeb_b_l[1:0]), .sp4_v_b(net294[0:15]),
     .sp4_h_l(sp4_v_b_01_00[47:0]), .sp12_h_l(sp12_v_b_01_00[23:0]),
     .prog(prog), .spi_ss_in_b(net502[0:1]),
     .tnl_op(bnl_op_01_00[7:0]), .lft_op(lft_op_01_00[7:0]),
     .bnl_op(lft_op_02_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[23:0]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_00[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_b_l), .fabric_out(net312));
io_col4_BOT_rev I_io_t02 ( .sdo(net313), .sdi(net278), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .sp4_v_t(net294[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_b_l[3:2]), .pado(pado_b_l[3:2]),
     .padeb(padeb_b_l[3:2]), .sp4_v_b(net329[0:15]),
     .sp4_h_l(sp4_v_b_02_00[47:0]), .sp12_h_l(sp12_v_b_02_00[23:0]),
     .prog(prog), .spi_ss_in_b(net333[0:1]),
     .tnl_op(lft_op_01_00[7:0]), .lft_op(lft_op_02_00[7:0]),
     .bnl_op(lft_op_03_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[47:24]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_00[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_b_l), .fabric_out(net494));
io_col4_BOT_rev I_io_t03 ( .sdo(net348), .sdi(net313), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .sp4_v_t(net329[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_b_l[5:4]), .pado(pado_b_l[5:4]),
     .padeb(padeb_b_l[5:4]), .sp4_v_b(net364[0:15]),
     .sp4_h_l(sp4_v_b_03_00[47:0]), .sp12_h_l(sp12_v_b_03_00[23:0]),
     .prog(prog), .spi_ss_in_b(net492[0:1]),
     .tnl_op(lft_op_02_00[7:0]), .lft_op(lft_op_03_00[7:0]),
     .bnl_op(lft_op_04_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[71:48]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_00[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_b_l), .fabric_out(net491));
io_col4_BOT_rev I_io_t05 ( .sdo(net383), .sdi(net418), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .sp4_v_t(net434[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_b_l[9:8]), .pado(pado_b_l[9:8]),
     .padeb(padeb_b_l[9:8]), .sp4_v_b(net399[0:15]),
     .sp4_h_l(sp4_v_b_05_00[47:0]), .sp12_h_l(sp12_v_b_05_00[23:0]),
     .prog(prog), .spi_ss_in_b(net497[0:1]),
     .tnl_op(lft_op_04_00[7:0]), .lft_op(lft_op_05_00[7:0]),
     .bnl_op(lft_op_06_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[119:96]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_00[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_b_l), .fabric_out(fabric_out_05_00));
io_col4_BOT_rev I_io_t04 ( .sdo(net418), .sdi(net348), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .sp4_v_t(net364[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_b_l[7:6]), .pado(pado_b_l[7:6]),
     .padeb(padeb_b_l[7:6]), .sp4_v_b(net434[0:15]),
     .sp4_h_l(sp4_v_b_04_00[47:0]), .sp12_h_l(sp12_v_b_04_00[23:0]),
     .prog(prog), .spi_ss_in_b(net501[0:1]),
     .tnl_op(lft_op_03_00[7:0]), .lft_op(lft_op_04_00[7:0]),
     .bnl_op(lft_op_05_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_04[5], bl_04[4], bl_04[37],
     bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32], bl_04[14],
     bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16], bl_04[27],
     bl_04[26], bl_04[25], bl_04[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[95:72]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_00[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_b_l), .fabric_out(net452));
io_col4_BOT_rev I_io_t06 ( .sdo(net453), .sdi(net383), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .sp4_v_t(net399[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_b_l[11:10]),
     .pado(pado_b_l[11:10]), .padeb(padeb_b_l[11:10]),
     .sp4_v_b(sp4_h_r_06_00[15:0]), .sp4_h_l(sp4_v_b_06_00[47:0]),
     .sp12_h_l(sp12_v_b_06_00[23:0]), .prog(prog),
     .spi_ss_in_b(net473[0:1]), .tnl_op(lft_op_05_00[7:0]),
     .lft_op(lft_op_06_00[7:0]), .bnl_op(tnr_op_06_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_06[5],
     bl_06[4], bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33],
     bl_06[32], bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17],
     bl_06[16], bl_06[27], bl_06[26], bl_06[25], bl_06[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_l[143:120]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_06_00[3:0]),
     .glb_netwk(glb_net_06[7:0]), .hold(hold_b_l),
     .fabric_out(fabric_out_06_00));
scanbuf1f I_scanbuf_mb ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(net453), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(tclk_o), .shift_o(shift_o),
     .sdo(sdo), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));

endmodule
// Library - leafcell, Cell - pinlatbuf12p, View - schematic
// LAST TIME SAVED: Mar 17 11:10:31 2009
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module pinlatbuf12p ( cout, cbit, icegate, pad_in, prog );
output  cout;

input  cbit, icegate, pad_in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I7 ( .A(net19), .Y(net024), .B(net13));
nand2_hvt I5 ( .A(icegate), .Y(net6), .B(cbit));
txgate_hvt I4 ( .in(cout), .out(net13), .pp(net6), .nn(net17));
txgate_hvt I1 ( .in(pad_in), .out(net13), .pp(net17), .nn(net6));
inv_hvt I6 ( .A(net6), .Y(net17));
inv_hvt I24 ( .A(prog), .Y(net19));
inv_hvt I23 ( .A(net024), .Y(cout));

endmodule
// Library - xpmem, Cell - cram2x2x6, View - schematic
// LAST TIME SAVED: Jul 28 08:29:06 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module cram2x2x6 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [23:0]  q;
output [23:0]  q_b;

inout [11:0]  bl;

input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  r_gnd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_5_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_base, View - schematic
// LAST TIME SAVED: Sep 13 06:51:33 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_base ( lc_trk_out, sp4_out, bl, min0, min1, min2,
     min3, pgate, prog, reset_b, sp12_in, vdd_cntl, wl );


input  prog;

output [1:0]  sp4_out;
output [3:0]  lc_trk_out;

inout [11:0]  bl;

input [1:0]  wl;
input [1:0]  sp12_in;
input [15:0]  min1;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [15:0]  min3;
input [1:0]  pgate;
input [15:0]  min0;
input [15:0]  min2;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  cbitb;

wire  [23:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
g_mux Imux2 ( .min(min2[15:0]), .prog(net60), .inmuxo(lc_trk_out[2]),
     .cbit({cbit[16], cbit[17], cbit[20], cbit[23], cbit[21]}),
     .cbitb({cbitb[16], cbitb[17], cbitb[20], cbitb[23], cbitb[21]}));
g_mux Imux3 ( .min(min3[15:0]), .prog(net60), .inmuxo(lc_trk_out[3]),
     .cbit({cbit[18], cbit[19], cbit[22], cbit[15], cbit[13]}),
     .cbitb({cbitb[18], cbitb[19], cbitb[22], cbitb[15], cbitb[13]}));
g_mux Imux1 ( .min(min1[15:0]), .prog(net60), .inmuxo(lc_trk_out[1]),
     .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}));
g_mux Imux0 ( .min(min0[15:0]), .prog(net60), .inmuxo(lc_trk_out[0]),
     .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}));
cram2x2x6 Imem2x2x6 ( .pgate(pgate[1:0]), .q(cbit[23:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[11:0]), .q_b(cbitb[23:0]));
sp12to4 Isp12to4_1_ ( .triout(sp4_out[1]), .cbitb(cbitb[11]),
     .drv(sp12_in[1]), .prog(net60));
sp12to4 Isp12to4_0_ ( .triout(sp4_out[0]), .cbitb(cbitb[9]),
     .drv(sp12_in[0]), .prog(net60));
inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net60));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0a, View - schematic
// LAST TIME SAVED: Jul 24 13:27:07 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_g0a ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g0;

inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;

input [7:0]  tnl_op;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  wl;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[34], sp4_r_v_b[25]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[33], sp4_r_v_b[26]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[35], sp4_r_v_b[24]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[32], sp4_r_v_b[27]}),
     .sp4_out(sp4_v_b[13:12]), .sp12_in({sp12_v_b[3], sp12_v_b[1]}),
     .lc_trk_out(lc_trk_g0[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0b, View - schematic
// LAST TIME SAVED: Jul 24 13:26:14 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_g0b ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, glb2local, lft_op,
     pgate, prog, reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op,
     vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g0;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
input [3:0]  glb2local;
input [7:0]  bnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  top_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], glb2local[1]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], glb2local[2]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], glb2local[0]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], glb2local[3]}),
     .sp4_out(sp4_v_b[15:14]), .sp12_in({sp12_v_b[7], sp12_v_b[5]}),
     .lc_trk_out(lc_trk_g0[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - xpmem, Cell - sg_bufx10, View - schematic
// LAST TIME SAVED: Jul 28 19:09:08 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module sg_bufx10 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1a, View - schematic
// LAST TIME SAVED: Jul 24 13:25:29 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_g1a ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [1:0]  wl;
input [7:0]  bnl_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[25], sp4_r_v_b[1]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[26], sp4_r_v_b[2]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[24], sp4_r_v_b[0]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[27], sp4_r_v_b[3]}),
     .sp4_out(sp4_v_b[17:16]), .sp12_in({sp12_v_b[11], sp12_v_b[9]}),
     .lc_trk_out(lc_trk_g1[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1b, View - schematic
// LAST TIME SAVED: Jul 24 13:24:39 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_g1b ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], sp4_r_v_b[5]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], sp4_r_v_b[6]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], sp4_r_v_b[4]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], sp4_r_v_b[7]}),
     .sp4_out(sp4_v_b[19:18]), .sp12_in({sp12_v_b[15], sp12_v_b[13]}),
     .lc_trk_out(lc_trk_g1[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2a, View - schematic
// LAST TIME SAVED: Jul 24 13:23:46 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_g2a ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g2;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;

input [7:0]  lft_op;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnl_op;
input [7:0]  slf_op;
input [1:0]  vdd_cntl;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  bnr_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[33], sp4_r_v_b[9]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[34], sp4_r_v_b[10]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[32], sp4_r_v_b[8]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[35], sp4_r_v_b[11]}),
     .sp4_out(sp4_v_b[21:20]), .sp12_in({sp12_v_b[19], sp12_v_b[17]}),
     .lc_trk_out(lc_trk_g2[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2b, View - schematic
// LAST TIME SAVED: Jul 24 13:22:58 2007
// NETLIST TIME: Aug 24 09:59:00 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_g2b ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g2;

inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [7:0]  bnr_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[37], sp4_r_v_b[13]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[38], sp4_r_v_b[14]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[36], sp4_r_v_b[12]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[39], sp4_r_v_b[15]}),
     .sp4_out(sp4_v_b[23:22]), .sp12_in({sp12_v_b[23], sp12_v_b[21]}),
     .lc_trk_out(lc_trk_g2[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3a, View - schematic
// LAST TIME SAVED: Jul 24 13:22:20 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_g3a ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g3;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  top_op;
input [1:0]  vdd_cntl;
input [7:0]  bnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  bnl_op;
input [7:0]  tnr_op;
input [7:0]  bot_op;
input [1:0]  wl;
input [7:0]  slf_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[41], sp4_r_v_b[17]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[42], sp4_r_v_b[18]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[40], sp4_r_v_b[16]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[43], sp4_r_v_b[19]}),
     .sp4_out(sp4_h_r[13:12]), .sp12_in({sp12_h_r[2], sp12_h_r[0]}),
     .lc_trk_out(lc_trk_g3[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3b, View - schematic
// LAST TIME SAVED: Jul 24 13:21:26 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module gmux_sp12to4_g3b ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g3;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;

input [7:0]  top_op;
input [7:0]  bnr_op;
input [1:0]  reset_b;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  wl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [1:0]  vdd_cntl;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[45], sp4_r_v_b[21]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[46], sp4_r_v_b[22]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[44], sp4_r_v_b[20]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[47], sp4_r_v_b[23]}),
     .sp4_out(sp4_h_r[15:14]), .sp12_in({sp12_h_r[6], sp12_h_r[4]}),
     .lc_trk_out(lc_trk_g3[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4, View - schematic
// LAST TIME SAVED: Jul 25 23:13:29 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module gmux_sp12to4 ( lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, bl,
     sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bnl_op, bnr_op,
     bot_op, glb2local, lft_op, pgate, prog, reset_b, rgt_op, slf_op,
     tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g3;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;

input [7:0]  slf_op;
input [7:0]  top_op;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [7:0]  bot_op;
input [7:0]  lft_op;
input [7:0]  tnl_op;
input [7:0]  bnr_op;
input [3:0]  glb2local;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  reset_b;
input [7:0]  bnl_op;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_g0a Ig0_30 ( .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp12_v_b(sp12_v_b[23:0]),
     .lc_trk_g0(lc_trk_g0[3:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[1:0]), .reset_b(reset_b[1:0]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g0b Ig0_74 ( .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]),
     .glb2local(glb2local[3:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .lc_trk_g0(lc_trk_g0[7:4]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[3:2]),
     .reset_b(reset_b[3:2]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g1a Ig1_30 ( .vdd_cntl(vdd_cntl[5:4]), .pgate(pgate[5:4]),
     .bl(bl[11:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]),
     .lft_op(lft_op[7:0]), .prog(prog), .rgt_op(rgt_op[7:0]),
     .reset_b(reset_b[5:4]), .slf_op(slf_op[7:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .wl(wl[5:4]), .lc_trk_g1(lc_trk_g1[3:0]));
gmux_sp12to4_g1b Ig1_74 ( .vdd_cntl(vdd_cntl[7:6]), .pgate(pgate[7:6]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .lc_trk_g1(lc_trk_g1[7:4]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[7:6]), .reset_b(reset_b[7:6]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g2a Ig2_30 ( .vdd_cntl(vdd_cntl[9:8]), .wl(wl[9:8]),
     .reset_b(reset_b[9:8]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[3:0]), .pgate(pgate[9:8]));
gmux_sp12to4_g2b Ig2_74 ( .vdd_cntl(vdd_cntl[11:10]),
     .pgate(pgate[11:10]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[11:10]),
     .reset_b(reset_b[11:10]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g3a Ig3_30 ( .vdd_cntl(vdd_cntl[13:12]), .wl(wl[13:12]),
     .reset_b(reset_b[13:12]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .pgate(pgate[13:12]), .lc_trk_g3(lc_trk_g3[3:0]));
gmux_sp12to4_g3b Ig3_74 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g3(lc_trk_g3[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .prog(prog),
     .bl(bl[11:0]), .reset_b(reset_b[15:14]), .wl(wl[15:14]));

endmodule
// Library - xpmem, Cell - cram2x2x5, View - schematic
// LAST TIME SAVED: Jul 28 08:25:47 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module cram2x2x5 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [19:0]  q_b;
output [19:0]  q;

inout [9:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  r_gnd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - sbox11to9_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:54:03 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox11to9_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[4]), .in5(t[10]), .in4(r[2]), .in3(r[10]),
     .in2(r[7]), .in1(b[10]), .in0(b[5]), .out(l[10]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[5]), .in5(t[11]), .in4(r[3]), .in3(r[11]),
     .in2(r[8]), .in1(b[11]), .in0(b[6]), .out(l[11]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[3]), .in5(t[9]), .in4(r[1]), .in3(r[9]),
     .in2(r[6]), .in1(b[9]), .in0(b[4]), .out(l[9]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[3]), .in5(r[9]), .in4(b[1]), .in3(b[9]),
     .in2(b[6]), .in1(l[9]), .in0(l[4]), .out(t[9]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[5]), .in5(r[11]), .in4(b[3]), .in3(b[11]),
     .in2(b[8]), .in1(l[11]), .in0(l[6]), .out(t[11]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[4]), .in5(r[10]), .in4(b[2]), .in3(b[10]),
     .in2(b[7]), .in1(l[10]), .in0(l[5]), .out(t[10]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox11to9_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:53:32 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox11to9_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  b;

input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[4]), .in5(b[10]), .in4(l[2]), .in3(l[10]),
     .in2(l[7]), .in1(t[10]), .in0(t[5]), .out(r[10]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[5]), .in5(b[11]), .in4(l[3]), .in3(l[11]),
     .in2(l[8]), .in1(t[11]), .in0(t[6]), .out(r[11]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[3]), .in5(b[9]), .in4(l[1]), .in3(l[9]),
     .in2(l[6]), .in1(t[9]), .in0(t[4]), .out(r[9]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[4]), .in5(l[10]), .in4(t[2]), .in3(t[10]),
     .in2(t[7]), .in1(r[10]), .in0(r[5]), .out(b[10]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[5]), .in5(l[11]), .in4(t[3]), .in3(t[11]),
     .in2(t[8]), .in1(r[11]), .in0(r[6]), .out(b[11]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[3]), .in5(l[9]), .in4(t[1]), .in3(t[9]),
     .in2(t[6]), .in1(r[9]), .in0(r[4]), .out(b[9]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - tiehi, View - schematic
// LAST TIME SAVED: Jul  8 16:18:10 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module tiehi ( tiehi );
output  tiehi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - leafcell, Cell - sbox8to6_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:52:49 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox8to6_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[1]), .in5(t[7]), .in4(r[11]), .in3(r[7]),
     .in2(r[4]), .in1(b[7]), .in0(b[2]), .out(l[7]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[2]), .in5(t[8]), .in4(r[0]), .in3(r[8]),
     .in2(r[5]), .in1(b[8]), .in0(b[3]), .out(l[8]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[0]), .in5(t[6]), .in4(r[10]), .in3(r[6]),
     .in2(r[3]), .in1(b[6]), .in0(b[1]), .out(l[6]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[0]), .in5(r[6]), .in4(b[10]), .in3(b[6]),
     .in2(b[3]), .in1(l[6]), .in0(l[1]), .out(t[6]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[2]), .in5(r[8]), .in4(b[0]), .in3(b[8]),
     .in2(b[5]), .in1(l[8]), .in0(l[3]), .out(t[8]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[1]), .in5(r[7]), .in4(b[11]), .in3(b[7]),
     .in2(b[4]), .in1(l[7]), .in0(l[2]), .out(t[7]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox8to6_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:36:51 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox8to6_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  cbit;

wire  [19:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[1]), .in5(b[7]), .in4(l[11]), .in3(l[7]),
     .in2(l[4]), .in1(t[7]), .in0(t[2]), .out(r[7]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[2]), .in5(b[8]), .in4(l[0]), .in3(l[8]),
     .in2(l[5]), .in1(t[8]), .in0(t[3]), .out(r[8]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[0]), .in5(b[6]), .in4(l[10]), .in3(l[6]),
     .in2(l[3]), .in1(t[6]), .in0(t[1]), .out(r[6]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[1]), .in5(l[7]), .in4(t[11]), .in3(t[7]),
     .in2(t[4]), .in1(r[7]), .in0(r[2]), .out(b[7]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[2]), .in5(l[8]), .in4(t[0]), .in3(t[8]),
     .in2(t[5]), .in1(r[8]), .in0(r[3]), .out(b[8]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[0]), .in5(l[6]), .in4(t[10]), .in3(t[6]),
     .in2(t[3]), .in1(r[6]), .in0(r[1]), .out(b[6]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox5to3_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:36:06 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox5to3_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  t;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[10]), .in5(t[4]), .in4(r[8]), .in3(r[4]),
     .in2(r[1]), .in1(b[4]), .in0(b[11]), .out(l[4]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[11]), .in5(t[5]), .in4(r[9]), .in3(r[5]),
     .in2(r[2]), .in1(b[5]), .in0(b[0]), .out(l[5]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[9]), .in5(t[3]), .in4(r[7]), .in3(r[3]),
     .in2(r[0]), .in1(b[3]), .in0(b[10]), .out(l[3]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[9]), .in5(r[3]), .in4(b[7]), .in3(b[3]),
     .in2(b[0]), .in1(l[3]), .in0(l[10]), .out(t[3]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[11]), .in5(r[5]), .in4(b[9]), .in3(b[5]),
     .in2(b[2]), .in1(l[5]), .in0(l[0]), .out(t[5]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[10]), .in5(r[4]), .in4(b[8]), .in3(b[4]),
     .in2(b[1]), .in1(l[4]), .in0(l[11]), .out(t[4]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 I534 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - sbox5to3_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:35:35 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox5to3_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;

input [1:0]  wl;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbitb;

wire  [19:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[10]), .in5(b[4]), .in4(l[8]), .in3(l[4]),
     .in2(l[1]), .in1(t[4]), .in0(t[11]), .out(r[4]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[11]), .in5(b[5]), .in4(l[9]), .in3(l[5]),
     .in2(l[2]), .in1(t[5]), .in0(t[0]), .out(r[5]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[9]), .in5(b[3]), .in4(l[7]), .in3(l[3]),
     .in2(l[0]), .in1(t[3]), .in0(t[10]), .out(r[3]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[10]), .in5(l[4]), .in4(t[8]), .in3(t[4]),
     .in2(t[1]), .in1(r[4]), .in0(r[11]), .out(b[4]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[11]), .in5(l[5]), .in4(t[9]), .in3(t[5]),
     .in2(t[2]), .in1(r[5]), .in0(r[0]), .out(b[5]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[9]), .in5(l[3]), .in4(t[7]), .in3(t[3]),
     .in2(t[0]), .in1(r[3]), .in0(r[10]), .out(b[3]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox2to0_220_p2, View - schematic
// LAST TIME SAVED: Nov 13 15:13:20 2008
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox2to0_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [11:0]  b;
inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  r;
inout [11:0]  l;

input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbitb;

wire  [19:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[7]), .in5(t[1]), .in4(r[5]), .in3(r[1]),
     .in2(r[10]), .in1(b[1]), .in0(b[8]), .out(l[1]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[8]), .in5(t[2]), .in4(r[6]), .in3(r[2]),
     .in2(r[11]), .in1(b[2]), .in0(b[9]), .out(l[2]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[6]), .in5(t[0]), .in4(r[4]), .in3(r[0]),
     .in2(r[9]), .in1(b[0]), .in0(b[7]), .out(l[0]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[6]), .in5(r[0]), .in4(b[4]), .in3(b[0]),
     .in2(b[9]), .in1(l[0]), .in0(l[7]), .out(t[0]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[8]), .in5(r[2]), .in4(b[6]), .in3(b[2]),
     .in2(b[11]), .in1(l[2]), .in0(l[9]), .out(t[2]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[7]), .in5(r[1]), .in4(b[5]), .in3(b[1]),
     .in2(b[10]), .in1(l[1]), .in0(l[8]), .out(t[1]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox2to0_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:34:25 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox2to0_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;
inout [9:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  cbit;

wire  [19:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[7]), .in5(b[1]), .in4(l[5]), .in3(l[1]),
     .in2(l[10]), .in1(t[1]), .in0(t[8]), .out(r[1]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[8]), .in5(b[2]), .in4(l[6]), .in3(l[2]),
     .in2(l[11]), .in1(t[2]), .in0(t[9]), .out(r[2]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[6]), .in5(b[0]), .in4(l[4]), .in3(l[0]),
     .in2(l[9]), .in1(t[0]), .in0(t[7]), .out(r[0]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[7]), .in5(l[1]), .in4(t[5]), .in3(t[1]),
     .in2(t[10]), .in1(r[1]), .in0(r[8]), .out(b[1]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[8]), .in5(l[2]), .in4(t[6]), .in3(t[2]),
     .in2(t[11]), .in1(r[2]), .in0(r[9]), .out(b[2]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[6]), .in5(l[0]), .in4(t[4]), .in3(t[0]),
     .in2(t[9]), .in1(r[0]), .in0(r[7]), .out(b[0]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - span4_switchandmem, View - schematic
// LAST TIME SAVED: Nov 13 15:13:23 2008
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module span4_switchandmem ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [11:0]  l;
inout [11:0]  t;
inout [11:0]  r;
inout [11:0]  b;
inout [9:0]  bl;

input [15:0]  vdd_cntl;
input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



sbox11to9_220_p2 I73 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .l(l[11:0]), .r(r[11:0]), .t(t[11:0]),
     .b(b[11:0]), .prog(prog), .wl(wl[15:14]), .bl(bl[9:0]),
     .reset_b(reset_b[15:14]));
sbox11to9_220_p1 I75 ( .vdd_cntl(vdd_cntl[13:12]),
     .pgate(pgate[13:12]), .l(l[11:0]), .r(r[11:0]), .t(t[11:0]),
     .b(b[11:0]), .prog(prog), .wl(wl[13:12]), .bl(bl[9:0]),
     .reset_b(reset_b[13:12]));
sbox8to6_220_p2 I74 ( .vdd_cntl(vdd_cntl[11:10]), .pgate(pgate[11:10]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[11:10]), .bl(bl[9:0]), .reset_b(reset_b[11:10]));
sbox8to6_220_p1 I76 ( .vdd_cntl(vdd_cntl[9:8]), .pgate(pgate[9:8]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[9:8]), .bl(bl[9:0]), .reset_b(reset_b[9:8]));
sbox5to3_220_p2 I71 ( .vdd_cntl(vdd_cntl[7:6]), .pgate(pgate[7:6]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[7:6]), .bl(bl[9:0]), .reset_b(reset_b[7:6]));
sbox5to3_220_p1 I72 ( .vdd_cntl(vdd_cntl[5:4]), .pgate(pgate[5:4]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[5:4]), .bl(bl[9:0]), .reset_b(reset_b[5:4]));
sbox2to0_220_p2 I70 ( .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[3:2]), .bl(bl[9:0]), .reset_b(reset_b[3:2]));
sbox2to0_220_p1 I69 ( .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[1:0]), .bl(bl[9:0]), .reset_b(reset_b[1:0]));

endmodule
// Library - leafcell, Cell - span4, View - schematic
// LAST TIME SAVED: Nov 13 15:13:26 2008
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module span4 ( bl, sp4_h_l, sp4_h_r, sp4_v_b, sp4_v_t, pgate, prog,
     reset_b, vdd_cntl, wl );

input  prog;

inout [47:0]  sp4_h_l;
inout [47:0]  sp4_h_r;
inout [9:0]  bl;
inout [47:0]  sp4_v_t;
inout [47:0]  sp4_v_b;

input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  wl;
input [15:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  sp4_h_r_mid;

wire  [11:0]  sp4_v_b_mid;



rm7  R1_27_ ( .MINUS(sp4_h_r[47]), .PLUS(sp4_h_l[34]));
rm7  R1_26_ ( .MINUS(sp4_h_r[46]), .PLUS(sp4_h_l[35]));
rm7  R1_25_ ( .MINUS(sp4_h_r[45]), .PLUS(sp4_h_l[32]));
rm7  R1_24_ ( .MINUS(sp4_h_r[44]), .PLUS(sp4_h_l[33]));
rm7  R1_23_ ( .MINUS(sp4_h_r[43]), .PLUS(sp4_h_l[30]));
rm7  R1_22_ ( .MINUS(sp4_h_r[42]), .PLUS(sp4_h_l[31]));
rm7  R1_21_ ( .MINUS(sp4_h_r[41]), .PLUS(sp4_h_l[28]));
rm7  R1_20_ ( .MINUS(sp4_h_r[40]), .PLUS(sp4_h_l[29]));
rm7  R1_19_ ( .MINUS(sp4_h_r[39]), .PLUS(sp4_h_l[26]));
rm7  R1_18_ ( .MINUS(sp4_h_r[38]), .PLUS(sp4_h_l[27]));
rm7  R1_17_ ( .MINUS(sp4_h_r[37]), .PLUS(sp4_h_l[24]));
rm7  R1_16_ ( .MINUS(sp4_h_r[36]), .PLUS(sp4_h_l[25]));
rm7  R1_15_ ( .MINUS(sp4_h_r[35]), .PLUS(sp4_h_l[22]));
rm7  R1_14_ ( .MINUS(sp4_h_r[34]), .PLUS(sp4_h_l[23]));
rm7  R1_13_ ( .MINUS(sp4_h_r[23]), .PLUS(sp4_h_l[10]));
rm7  R1_12_ ( .MINUS(sp4_h_r[22]), .PLUS(sp4_h_l[11]));
rm7  R1_11_ ( .MINUS(sp4_h_r_mid[11]), .PLUS(sp4_h_l[46]));
rm7  R1_10_ ( .MINUS(sp4_h_r_mid[10]), .PLUS(sp4_h_l[47]));
rm7  R1_9_ ( .MINUS(sp4_h_r_mid[9]), .PLUS(sp4_h_l[44]));
rm7  R1_8_ ( .MINUS(sp4_h_r_mid[8]), .PLUS(sp4_h_l[45]));
rm7  R1_7_ ( .MINUS(sp4_h_r_mid[7]), .PLUS(sp4_h_l[42]));
rm7  R1_6_ ( .MINUS(sp4_h_r_mid[6]), .PLUS(sp4_h_l[43]));
rm7  R1_5_ ( .MINUS(sp4_h_r_mid[5]), .PLUS(sp4_h_l[40]));
rm7  R1_4_ ( .MINUS(sp4_h_r_mid[4]), .PLUS(sp4_h_l[41]));
rm7  R1_3_ ( .MINUS(sp4_h_r_mid[3]), .PLUS(sp4_h_l[38]));
rm7  R1_2_ ( .MINUS(sp4_h_r_mid[2]), .PLUS(sp4_h_l[39]));
rm7  R1_1_ ( .MINUS(sp4_h_r_mid[1]), .PLUS(sp4_h_l[36]));
rm7  R1_0_ ( .MINUS(sp4_h_r_mid[0]), .PLUS(sp4_h_l[37]));
rm5  R2_19_ ( .MINUS(sp4_h_r[33]), .PLUS(sp4_h_l[20]));
rm5  R2_18_ ( .MINUS(sp4_h_r[32]), .PLUS(sp4_h_l[21]));
rm5  R2_17_ ( .MINUS(sp4_h_r[31]), .PLUS(sp4_h_l[18]));
rm5  R2_16_ ( .MINUS(sp4_h_r[30]), .PLUS(sp4_h_l[19]));
rm5  R2_15_ ( .MINUS(sp4_h_r[29]), .PLUS(sp4_h_l[16]));
rm5  R2_14_ ( .MINUS(sp4_h_r[28]), .PLUS(sp4_h_l[17]));
rm5  R2_13_ ( .MINUS(sp4_h_r[27]), .PLUS(sp4_h_l[14]));
rm5  R2_12_ ( .MINUS(sp4_h_r[26]), .PLUS(sp4_h_l[15]));
rm5  R2_11_ ( .MINUS(sp4_h_r[25]), .PLUS(sp4_h_l[12]));
rm5  R2_10_ ( .MINUS(sp4_h_r[24]), .PLUS(sp4_h_l[13]));
rm5  R2_9_ ( .MINUS(sp4_h_r[21]), .PLUS(sp4_h_l[8]));
rm5  R2_8_ ( .MINUS(sp4_h_r[20]), .PLUS(sp4_h_l[9]));
rm5  R2_7_ ( .MINUS(sp4_h_r[19]), .PLUS(sp4_h_l[6]));
rm5  R2_6_ ( .MINUS(sp4_h_r[18]), .PLUS(sp4_h_l[7]));
rm5  R2_5_ ( .MINUS(sp4_h_r[17]), .PLUS(sp4_h_l[4]));
rm5  R2_4_ ( .MINUS(sp4_h_r[16]), .PLUS(sp4_h_l[5]));
rm5  R2_3_ ( .MINUS(sp4_h_r[15]), .PLUS(sp4_h_l[2]));
rm5  R2_2_ ( .MINUS(sp4_h_r[14]), .PLUS(sp4_h_l[3]));
rm5  R2_1_ ( .MINUS(sp4_h_r[13]), .PLUS(sp4_h_l[0]));
rm5  R2_0_ ( .MINUS(sp4_h_r[12]), .PLUS(sp4_h_l[1]));
rm6  R0_47_ ( .MINUS(sp4_v_b[47]), .PLUS(sp4_v_t[34]));
rm6  R0_46_ ( .MINUS(sp4_v_b[46]), .PLUS(sp4_v_t[35]));
rm6  R0_45_ ( .MINUS(sp4_v_b[45]), .PLUS(sp4_v_t[32]));
rm6  R0_44_ ( .MINUS(sp4_v_b[44]), .PLUS(sp4_v_t[33]));
rm6  R0_43_ ( .MINUS(sp4_v_b[43]), .PLUS(sp4_v_t[30]));
rm6  R0_42_ ( .MINUS(sp4_v_b[42]), .PLUS(sp4_v_t[31]));
rm6  R0_41_ ( .MINUS(sp4_v_b[41]), .PLUS(sp4_v_t[28]));
rm6  R0_40_ ( .MINUS(sp4_v_b[40]), .PLUS(sp4_v_t[29]));
rm6  R0_39_ ( .MINUS(sp4_v_b[39]), .PLUS(sp4_v_t[26]));
rm6  R0_38_ ( .MINUS(sp4_v_b[38]), .PLUS(sp4_v_t[27]));
rm6  R0_37_ ( .MINUS(sp4_v_b[37]), .PLUS(sp4_v_t[24]));
rm6  R0_36_ ( .MINUS(sp4_v_b[36]), .PLUS(sp4_v_t[25]));
rm6  R0_35_ ( .MINUS(sp4_v_b[35]), .PLUS(sp4_v_t[22]));
rm6  R0_34_ ( .MINUS(sp4_v_b[34]), .PLUS(sp4_v_t[23]));
rm6  R0_33_ ( .MINUS(sp4_v_b[33]), .PLUS(sp4_v_t[20]));
rm6  R0_32_ ( .MINUS(sp4_v_b[32]), .PLUS(sp4_v_t[21]));
rm6  R0_31_ ( .MINUS(sp4_v_b[31]), .PLUS(sp4_v_t[18]));
rm6  R0_30_ ( .MINUS(sp4_v_b[30]), .PLUS(sp4_v_t[19]));
rm6  R0_29_ ( .MINUS(sp4_v_b[29]), .PLUS(sp4_v_t[16]));
rm6  R0_28_ ( .MINUS(sp4_v_b[28]), .PLUS(sp4_v_t[17]));
rm6  R0_27_ ( .MINUS(sp4_v_b[27]), .PLUS(sp4_v_t[14]));
rm6  R0_26_ ( .MINUS(sp4_v_b[26]), .PLUS(sp4_v_t[15]));
rm6  R0_25_ ( .MINUS(sp4_v_b[25]), .PLUS(sp4_v_t[12]));
rm6  R0_24_ ( .MINUS(sp4_v_b[24]), .PLUS(sp4_v_t[13]));
rm6  R0_23_ ( .MINUS(sp4_v_b[23]), .PLUS(sp4_v_t[10]));
rm6  R0_22_ ( .MINUS(sp4_v_b[22]), .PLUS(sp4_v_t[11]));
rm6  R0_21_ ( .MINUS(sp4_v_b[21]), .PLUS(sp4_v_t[8]));
rm6  R0_20_ ( .MINUS(sp4_v_b[20]), .PLUS(sp4_v_t[9]));
rm6  R0_19_ ( .MINUS(sp4_v_b[19]), .PLUS(sp4_v_t[6]));
rm6  R0_18_ ( .MINUS(sp4_v_b[18]), .PLUS(sp4_v_t[7]));
rm6  R0_17_ ( .MINUS(sp4_v_b[17]), .PLUS(sp4_v_t[4]));
rm6  R0_16_ ( .MINUS(sp4_v_b[16]), .PLUS(sp4_v_t[5]));
rm6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[2]));
rm6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[3]));
rm6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[0]));
rm6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[1]));
rm6  R0_11_ ( .MINUS(sp4_v_b_mid[11]), .PLUS(sp4_v_t[46]));
rm6  R0_10_ ( .MINUS(sp4_v_b_mid[10]), .PLUS(sp4_v_t[47]));
rm6  R0_9_ ( .MINUS(sp4_v_b_mid[9]), .PLUS(sp4_v_t[44]));
rm6  R0_8_ ( .MINUS(sp4_v_b_mid[8]), .PLUS(sp4_v_t[45]));
rm6  R0_7_ ( .MINUS(sp4_v_b_mid[7]), .PLUS(sp4_v_t[42]));
rm6  R0_6_ ( .MINUS(sp4_v_b_mid[6]), .PLUS(sp4_v_t[43]));
rm6  R0_5_ ( .MINUS(sp4_v_b_mid[5]), .PLUS(sp4_v_t[40]));
rm6  R0_4_ ( .MINUS(sp4_v_b_mid[4]), .PLUS(sp4_v_t[41]));
rm6  R0_3_ ( .MINUS(sp4_v_b_mid[3]), .PLUS(sp4_v_t[38]));
rm6  R0_2_ ( .MINUS(sp4_v_b_mid[2]), .PLUS(sp4_v_t[39]));
rm6  R0_1_ ( .MINUS(sp4_v_b_mid[1]), .PLUS(sp4_v_t[36]));
rm6  R0_0_ ( .MINUS(sp4_v_b_mid[0]), .PLUS(sp4_v_t[37]));
span4_switchandmem ISPAN4_SW ( .vdd_cntl(vdd_cntl[15:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]), .b(sp4_v_b[11:0]),
     .r(sp4_h_r[11:0]), .l(sp4_h_r_mid[11:0]), .prog(prog),
     .wl(wl[15:0]), .t(sp4_v_b_mid[11:0]), .bl(bl[9:0]));

endmodule
// Library - leafcell, Cell - clkmandcmuxrev0, View - schematic
// LAST TIME SAVED: Nov 14 11:27:18 2008
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module clkmandcmuxrev0 ( clk, clkb, glb2local, s_r, cbit, cbitb,
     glb_netwk, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, min0, min1,
     min2, min3, prog );
output  clk, clkb, s_r;

input  prog;

output [3:0]  glb2local;

input [7:0]  min1;
input [7:0]  min3;
input [7:0]  min2;
input [31:0]  cbitb;
input [7:0]  min0;
input [31:0]  cbit;
input [7:0]  glb_netwk;
input [5:0]  lc_trk_g0;
input [5:0]  lc_trk_g1;
input [5:0]  lc_trk_g2;
input [5:0]  lc_trk_g3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



sr_clkm8to1 I_srmux8to1 ( .mout(s_r), .cbitb(cbitb[12:9]),
     .min({lc_trk_g3[5], lc_trk_g2[4], lc_trk_g1[5], lc_trk_g0[4],
     glb_netwk[6], glb_netwk[4], glb_netwk[2], glb_netwk[0]}),
     .cbit(cbit[12:9]), .prog(prog));
ce_clkm8to1 I_cemux8to1 ( .cbitb(cbitb[8:5]), .min({lc_trk_g3[3],
     lc_trk_g2[2], lc_trk_g1[3], lc_trk_g0[2], glb_netwk[7],
     glb_netwk[5], glb_netwk[3], glb_netwk[1]}), .cbit(cbit[8:5]),
     .moutb(ceb), .prog(prog));
clk_mux12to1 I_clkmux12to1 ( .min({lc_trk_g3[1], lc_trk_g2[0],
     lc_trk_g1[1], lc_trk_g0[0], glb_netwk[7:0]}), .clk(clk),
     .clkb(clkb), .cbitb({cbitb[31], cbitb[4], cbitb[3], cbitb[2],
     cbitb[1], cbitb[0]}), .cbit({cbit[31], cbit[4], cbit[3], cbit[2],
     cbit[1], cbit[0]}), .cenb(ceb), .prog(prog));
clk_mux8to1 I_clkmux8to1_1 ( .prog(prog), .inmuxo(glb2local[1]),
     .min(min2[7:0]), .cbit(cbit[20:17]), .cbitb(cbitb[20:17]));
clk_mux8to1 I_clkmux8to1_2 ( .prog(prog), .inmuxo(glb2local[2]),
     .min(min1[7:0]), .cbit(cbit[24:21]), .cbitb(cbitb[24:21]));
clk_mux8to1 I_clkmux8to1_3 ( .prog(prog), .inmuxo(glb2local[3]),
     .min(min0[7:0]), .cbit(cbit[28:25]), .cbitb(cbitb[28:25]));
clk_mux8to1 I_clkmux8to1_0 ( .inmuxo(glb2local[0]), .min(min3[7:0]),
     .cbit(cbit[16:13]), .cbitb(cbitb[16:13]), .prog(prog));

endmodule
// Library - leafcell, Cell - sbox1, View - schematic
// LAST TIME SAVED: Nov 13 16:05:04 2008
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module sbox1 ( b, l, r, t, c, cb, prog );
inout  b, l, r, t;

input  prog;

input [7:0]  c;
input [7:0]  cb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



sbox1m3to1 I232 ( .in2(r), .cb(cb[7:6]), .op(t), .in0(l), .in1(b),
     .c(c[7:6]), .prog(prog));
sbox1m3to1 I230 ( .in2(r), .cb(cb[3:2]), .op(l), .in0(b), .in1(t),
     .c(c[3:2]), .prog(prog));
sbox1m3to1 I226 ( .in2(r), .cb(cb[1:0]), .op(b), .in0(l), .in1(t),
     .c(c[1:0]), .prog(prog));
sbox1m3to1 I231 ( .in2(b), .cb(cb[5:4]), .op(r), .in0(l), .in1(t),
     .c(c[5:4]), .prog(prog));

endmodule
// Library - misc, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jul  3 16:54:18 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_dff ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));
nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));

endmodule
// Library - xpmem, Cell - cram16x4, View - schematic
// LAST TIME SAVED: Jul 28 08:31:30 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module cram16x4 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [63:0]  q_b;
output [63:0]  q;

inout [3:0]  bl;

input [15:0]  pgate;
input [15:0]  r_gnd;
input [15:0]  wl;
input [15:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 I16_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[1:0]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[15:14]));
cram2x2 I16_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[1:0]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[13:12]));
cram2x2 I16_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[1:0]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[11:10]));
cram2x2 I16_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[1:0]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[9:8]));
cram2x2 I16_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[1:0]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[7:6]));
cram2x2 I16_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[1:0]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[5:4]));
cram2x2 I16_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[1:0]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[3:2]));
cram2x2 I16_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[3:2]), .q_b(q_b[63:60]),
     .q(q[63:60]), .wl(wl[15:14]));
cram2x2 Imstake_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[3:2]), .q_b(q_b[59:56]),
     .q(q[59:56]), .wl(wl[13:12]));
cram2x2 Imstake_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[3:2]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[11:10]));
cram2x2 Imstake_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[3:2]), .q_b(q_b[51:48]), .q(q[51:48]),
     .wl(wl[9:8]));
cram2x2 Imstake_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[3:2]), .q_b(q_b[47:44]), .q(q[47:44]),
     .wl(wl[7:6]));
cram2x2 Imstake_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[3:2]), .q_b(q_b[43:40]), .q(q[43:40]),
     .wl(wl[5:4]));
cram2x2 Imstake_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[3:2]), .q_b(q_b[39:36]), .q(q[39:36]),
     .wl(wl[3:2]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[35:32]), .q(q[35:32]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - misc_module4rev0, View - schematic
// LAST TIME SAVED: Jan 20 08:53:58 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module misc_module4rev0 ( S_R, .cbit_colcntl({cbit[60], cbit[56],
     cbit[52], cbit[48], cbit[44], cbit[40], cbit[32], cbit[3]}), clk,
     clkb, glb2local, sp4, bl, b, glb_netwk, l, lc_trk_g0, lc_trk_g1,
     lc_trk_g2, lc_trk_g3, m, min0, min1, min2, min3, pgate, prog, r,
     reset_b, sp12, vdd_cntl, wl );
output  S_R, clk, clkb;


input  prog;

output [7:0]  sp4;
output [3:0]  glb2local;
output [63:0]  cbit;

inout [3:0]  bl;

input [7:0]  sp12;
input [5:0]  lc_trk_g3;
input [15:0]  wl;
input [5:0]  lc_trk_g1;
input [1:0]  b;
input [15:0]  vdd_cntl;
input [1:0]  r;
input [7:0]  min3;
input [15:0]  pgate;
input [5:0]  lc_trk_g0;
input [7:0]  glb_netwk;
input [7:0]  min1;
input [1:0]  m;
input [7:0]  min0;
input [7:0]  min2;
input [15:0]  reset_b;
input [5:0]  lc_trk_g2;
input [1:0]  l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  r_vdd;

wire  [63:0]  cbitb;



clkmandcmuxrev0 I_tclkmux ( .prog(prog), .min3(min3[7:0]),
     .min2(min2[7:0]), .min1(min1[7:0]), .min0(min0[7:0]),
     .lc_trk_g3(lc_trk_g3[5:0]), .lc_trk_g2(lc_trk_g2[5:0]),
     .lc_trk_g1(lc_trk_g1[5:0]), .lc_trk_g0(lc_trk_g0[5:0]),
     .glb_netwk(glb_netwk[7:0]), .cbitb({cbitb[2], cbitb[1], cbitb[0],
     cbitb[27], cbitb[25], cbitb[26], cbitb[24], cbitb[23], cbitb[21],
     cbitb[22], cbitb[20], cbitb[19], cbitb[17], cbitb[18], cbitb[16],
     cbitb[15], cbitb[13], cbitb[14], cbitb[12], cbitb[31], cbitb[29],
     cbitb[30], cbitb[28], cbitb[11], cbitb[9], cbitb[10], cbitb[8],
     cbitb[38], cbitb[36], cbitb[7], cbitb[6], cbitb[4]}),
     .cbit({cbit[2], cbit[1], cbit[0], cbit[27], cbit[25], cbit[26],
     cbit[24], cbit[23], cbit[21], cbit[22], cbit[20], cbit[19],
     cbit[17], cbit[18], cbit[16], cbit[15], cbit[13], cbit[14],
     cbit[12], cbit[31], cbit[29], cbit[30], cbit[28], cbit[11],
     cbit[9], cbit[10], cbit[8], cbit[38], cbit[36], cbit[7], cbit[6],
     cbit[4]}), .s_r(S_R), .glb2local(glb2local[3:0]), .clkb(clkb),
     .clk(clk));
pch_hvt  vdd_cntrl_15_ ( .D(r_vdd[15]), .B(vdd_), .G(vdd_cntl[15]),
     .S(vdd_));
pch_hvt  vdd_cntrl_14_ ( .D(r_vdd[14]), .B(vdd_), .G(vdd_cntl[14]),
     .S(vdd_));
pch_hvt  vdd_cntrl_13_ ( .D(r_vdd[13]), .B(vdd_), .G(vdd_cntl[13]),
     .S(vdd_));
pch_hvt  vdd_cntrl_12_ ( .D(r_vdd[12]), .B(vdd_), .G(vdd_cntl[12]),
     .S(vdd_));
pch_hvt  vdd_cntrl_11_ ( .D(r_vdd[11]), .B(vdd_), .G(vdd_cntl[11]),
     .S(vdd_));
pch_hvt  vdd_cntrl_10_ ( .D(r_vdd[10]), .B(vdd_), .G(vdd_cntl[10]),
     .S(vdd_));
pch_hvt  vdd_cntrl_9_ ( .D(r_vdd[9]), .B(vdd_), .G(vdd_cntl[9]),
     .S(vdd_));
pch_hvt  vdd_cntrl_8_ ( .D(r_vdd[8]), .B(vdd_), .G(vdd_cntl[8]),
     .S(vdd_));
pch_hvt  vdd_cntrl_7_ ( .D(r_vdd[7]), .B(vdd_), .G(vdd_cntl[7]),
     .S(vdd_));
pch_hvt  vdd_cntrl_6_ ( .D(r_vdd[6]), .B(vdd_), .G(vdd_cntl[6]),
     .S(vdd_));
pch_hvt  vdd_cntrl_5_ ( .D(r_vdd[5]), .B(vdd_), .G(vdd_cntl[5]),
     .S(vdd_));
pch_hvt  vdd_cntrl_4_ ( .D(r_vdd[4]), .B(vdd_), .G(vdd_cntl[4]),
     .S(vdd_));
pch_hvt  vdd_cntrl_3_ ( .D(r_vdd[3]), .B(vdd_), .G(vdd_cntl[3]),
     .S(vdd_));
pch_hvt  vdd_cntrl_2_ ( .D(r_vdd[2]), .B(vdd_), .G(vdd_cntl[2]),
     .S(vdd_));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sp12to4 I_sp12to4_7_ ( .prog(progd), .triout(sp4[7]),
     .cbitb(cbitb[62]), .drv(sp12[7]));
sp12to4 I_sp12to4_6_ ( .prog(progd), .triout(sp4[6]),
     .cbitb(cbitb[58]), .drv(sp12[6]));
sp12to4 I_sp12to4_5_ ( .prog(progd), .triout(sp4[5]),
     .cbitb(cbitb[54]), .drv(sp12[5]));
sp12to4 I_sp12to4_4_ ( .prog(progd), .triout(sp4[4]),
     .cbitb(cbitb[50]), .drv(sp12[4]));
sp12to4 I_sp12to4_3_ ( .prog(progd), .triout(sp4[3]),
     .cbitb(cbitb[46]), .drv(sp12[3]));
sp12to4 I_sp12to4_2_ ( .prog(progd), .triout(sp4[2]),
     .cbitb(cbitb[42]), .drv(sp12[2]));
sp12to4 I_sp12to4_1_ ( .prog(progd), .triout(sp4[1]), .cbitb(cbitb[5]),
     .drv(sp12[1]));
sp12to4 I_sp12to4_0_ ( .prog(progd), .triout(sp4[0]),
     .cbitb(cbitb[34]), .drv(sp12[0]));
sbox1 I_span12_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(prog));
sbox1 I_span12_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(prog));
cram16x4 Ic64 ( .r_gnd(r_vdd[15:0]), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .q(cbit[63:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));
inv_hvt I76 ( .A(prog), .Y(progb));
inv_hvt I75 ( .A(progb), .Y(progd));

endmodule
// Library - leafcell, Cell - logic_cell, View - schematic
// LAST TIME SAVED: Aug 28 17:23:08 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module logic_cell ( carry_out, out, carry_in, cbit, clk, clkb, in0,
     in1, in2, in3, prog, purst, s_r );
output  carry_out, out;

input  carry_in, clk, clkb, in0, in1, in2, in3, prog, purst, s_r;

input [20:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



coredffr REG ( .purst(purst), .d(LUT4_outd), .q(rego),
     .cbit(cbit[17:16]), .clkb(clkb), .clk(clk), .S_R(s_r));
carry_logic ICARRY_LOGIC ( .b_bar(in1b1), .carry_in(carry_in), .b(in1),
     .cout(carry_out), .a(in2), .a_bar(in2b1), .vg_en(cbit[20]));
o_mux Iomux ( .in1(rego), .out(out), .cbit(cbit[19]), .prog(prog),
     .in0(LUT4_outd));
clut4 iclut4 ( .in0b(in0b1), .in3b(in3b1), .in2b(in2b1),
     .lut4(LUT4_outd), .in1b(in1b1), .in2(in2), .in1(in1), .in0(in0),
     .in3(in3), .cbit(cbit[15:0]));
inv_hvt I163 ( .A(in3), .Y(in3b1));
inv_hvt I164 ( .A(in1), .Y(in1b1));
inv_hvt I162 ( .A(in2), .Y(in2b1));
inv_hvt I161 ( .A(in0), .Y(in0b1));

endmodule
// Library - leafcell, Cell - odrv12_30, View - schematic
// LAST TIME SAVED: Jun  5 15:34:53 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module odrv12_30 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_h_r;

input  prog, slfop;

output [2:0]  sp4_h_r;
output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_r_v_b;

input [11:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



odrv12 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b[1]));
odrv12 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp12(sp12_v_b[0]));
odrv12 I70 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r));
odrv4 I69_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I71_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[2]));
odrv4 I71_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[1]));
odrv4 I71_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp4(sp4_v_b[0]));
odrv4 I73_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I73_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I73_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - xpmem, Cell - cram_2x28, View - schematic
// LAST TIME SAVED: Jul 28 08:32:33 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module cram_2x28 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [55:0]  q;
output [55:0]  q_b;

inout [27:0]  bl;

input [1:0]  wl;
input [1:0]  reset;
input [1:0]  r_vdd;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_13_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[27:26]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[1:0]));
cram2x2 Imstake_12_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[25:24]), .q_b(q_b[51:48]),
     .q(q[51:48]), .wl(wl[1:0]));
cram2x2 Imstake_11_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[23:22]), .q_b(q_b[47:44]),
     .q(q[47:44]), .wl(wl[1:0]));
cram2x2 Imstake_10_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[21:20]), .q_b(q_b[43:40]),
     .q(q[43:40]), .wl(wl[1:0]));
cram2x2 Imstake_9_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[19:18]), .q_b(q_b[39:36]),
     .q(q[39:36]), .wl(wl[1:0]));
cram2x2 Imstake_8_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[17:16]), .q_b(q_b[35:32]),
     .q(q[35:32]), .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[15:14]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[1:0]));
cram2x2 Imstake_6_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[13:12]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[1:0]));
cram2x2 Imstake_5_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - lcmuxod3_0rev, View - schematic
// LAST TIME SAVED: Jun  2 13:13:15 2008
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module lcmuxod3_0rev ( carry_out, cbit, cbitb, op, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1,
     min2, min3, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, sp12_h_r;

input  carry_in, clk, clkb, prog, purst, s_r;

output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;
output [55:0]  cbit;
output [55:0]  cbitb;

input [15:0]  min3;
input [27:0]  bl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [15:0]  min2;
input [15:0]  min0;
input [1:0]  reset_b;
input [1:0]  wl;
input [15:0]  min1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
logic_cell ILC ( .purst(purst), .in1(in1), .in3(in3), .in2(in2),
     .in0(in0), .s_r(s_r), .cbit({cbit[38], cbit[39], cbit[39],
     cbit[37], cbit[36], cbit[22], cbit[20], cbit[21], cbit[23],
     cbit[26], cbit[24], cbit[25], cbit[27], cbit[35], cbit[33],
     cbit[32], cbit[34], cbit[31], cbit[29], cbit[28], cbit[30]}),
     .prog(prog), .clkb(clkb), .carry_in(carry_in),
     .carry_out(carry_out), .clk(clk), .out(op));
in_mux in1mux ( .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}),
     .min(min1[15:0]), .prog(prog), .inmuxo(in1));
in_mux in0mux ( .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}),
     .min(min0[15:0]), .prog(prog), .inmuxo(in0));
in_mux in2mux ( .cbit({cbit[12], cbit[13], cbit[16], cbit[19],
     cbit[17]}), .cbitb({cbitb[12], cbitb[13], cbitb[16], cbitb[19],
     cbitb[17]}), .min(min2[15:0]), .prog(prog), .inmuxo(in2));
in_mux in3mux ( .min(min3[15:0]), .cbit({cbit[14], cbit[15], cbit[18],
     cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15], cbitb[18],
     cbitb[11], cbitb[9]}), .prog(prog), .inmuxo(in3));
odrv12_30 Iodrv30 ( .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53],
     cbitb[55], cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44],
     cbitb[46], cbitb[43], cbitb[41], cbitb[42], cbitb[40]}),
     .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_h_r(sp4_h_r[2:0]), .slfop(op),
     .prog(prog));
cram_2x28 I41 ( .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]), .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .q_b(cbitb[55:0]));

endmodule
// Library - leafcell, Cell - lcmuxod3_0, View - schematic
// LAST TIME SAVED: Aug 21 17:57:09 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module lcmuxod3_0 ( carry_out, op, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, sp12_h_r;

input  carry_in, clk, clkb, prog, purst, s_r;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_v_b;
output [2:0]  sp4_v_b;

input [15:0]  min2;
input [1:0]  wl;
input [15:0]  min3;
input [15:0]  min0;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [27:0]  bl;
input [1:0]  pgate;
input [15:0]  min1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
logic_cell ILC ( .purst(purst), .in1(in1), .in3(in3), .in2(in2),
     .in0(in0), .s_r(s_r), .cbit({cbit[38], cbit[39], cbit[39],
     cbit[37], cbit[36], cbit[22], cbit[20], cbit[21], cbit[23],
     cbit[26], cbit[24], cbit[25], cbit[27], cbit[35], cbit[33],
     cbit[32], cbit[34], cbit[31], cbit[29], cbit[28], cbit[30]}),
     .prog(prog), .clkb(clkb), .carry_in(carry_in),
     .carry_out(carry_out), .clk(clk), .out(op));
in_mux in1mux ( .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}),
     .min(min1[15:0]), .prog(prog), .inmuxo(in1));
in_mux in0mux ( .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}),
     .min(min0[15:0]), .prog(prog), .inmuxo(in0));
in_mux in2mux ( .cbit({cbit[12], cbit[13], cbit[16], cbit[19],
     cbit[17]}), .cbitb({cbitb[12], cbitb[13], cbitb[16], cbitb[19],
     cbitb[17]}), .min(min2[15:0]), .prog(prog), .inmuxo(in2));
in_mux in3mux ( .min(min3[15:0]), .cbit({cbit[14], cbit[15], cbit[18],
     cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15], cbitb[18],
     cbitb[11], cbitb[9]}), .prog(prog), .inmuxo(in3));
odrv12_30 Iodrv30 ( .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53],
     cbitb[55], cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44],
     cbitb[46], cbitb[43], cbitb[41], cbitb[42], cbitb[40]}),
     .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_h_r(sp4_h_r[2:0]), .slfop(op),
     .prog(prog));
cram_2x28 I41 ( .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]), .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .q_b(cbitb[55:0]));

endmodule
// Library - leafcell, Cell - odrv12_74, View - schematic
// LAST TIME SAVED: Jun  5 15:30:49 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module odrv12_74 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_v_b;

input  prog, slfop;

output [2:0]  sp4_v_b;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_h_r;

input [11:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



odrv12 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp12(sp12_h_r[1]));
odrv12 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r[0]));
odrv12 I71 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b));
odrv4 I68_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I68_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I68_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I70_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp4(sp4_v_b[2]));
odrv4 I70_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[1]));
odrv4 I70_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[0]));
odrv4 I72_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - lcmuxod7_4, View - schematic
// LAST TIME SAVED: Aug 21 17:56:42 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module lcmuxod7_4 ( carry_out, op, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, sp12_v_b;

input  carry_in, clk, clkb, prog, purst, s_r;

output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;
output [1:0]  sp12_h_r;
output [2:0]  sp4_v_b;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [15:0]  min2;
input [1:0]  reset_b;
input [15:0]  min3;
input [15:0]  min0;
input [27:0]  bl;
input [15:0]  min1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
in_mux in1mux ( .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}),
     .min(min1[15:0]), .prog(prog), .inmuxo(in1));
in_mux in0mux ( .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}),
     .min(min0[15:0]), .prog(prog), .inmuxo(in0));
in_mux in2mux ( .cbit({cbit[12], cbit[13], cbit[16], cbit[19],
     cbit[17]}), .cbitb({cbitb[12], cbitb[13], cbitb[16], cbitb[19],
     cbitb[17]}), .min(min2[15:0]), .prog(prog), .inmuxo(in2));
in_mux in3mux ( .min(min3[15:0]), .cbit({cbit[14], cbit[15], cbit[18],
     cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15], cbitb[18],
     cbitb[11], cbitb[9]}), .prog(prog), .inmuxo(in3));
logic_cell ILC ( .purst(purst), .in1(in1), .in3(in3), .in2(in2),
     .in0(in0), .s_r(s_r), .cbit({cbit[38], cbit[39], cbit[39],
     cbit[37], cbit[36], cbit[22], cbit[20], cbit[21], cbit[23],
     cbit[26], cbit[24], cbit[25], cbit[27], cbit[35], cbit[33],
     cbit[32], cbit[34], cbit[31], cbit[29], cbit[28], cbit[30]}),
     .prog(prog), .clkb(clkb), .carry_in(carry_in),
     .carry_out(carry_out), .clk(clk), .out(op));
odrv12_74 Iodrv74 ( .cbitb({cbitb[53], cbitb[55], cbitb[52], cbitb[54],
     cbitb[51], cbitb[49], cbitb[44], cbitb[46], cbitb[43], cbitb[41],
     cbitb[42], cbitb[40]}), .sp4_r_v_b(sp4_r_v_b[2:0]),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_h_r(sp4_h_r[2:0]),
     .sp12_v_b(sp12_v_b), .sp12_h_r(sp12_h_r[1:0]), .slfop(op),
     .prog(prog));
cram_2x28 I41 ( .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]), .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .q_b(cbitb[55:0]));

endmodule
// Library - leafcell, Cell - lccol_rev0, View - schematic
// LAST TIME SAVED: Jan 20 09:55:16 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module lccol_rev0 ( carry_out, slf_op, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, cin2local, clk, clkb, lc_trk_g0, lc_trk_g1,
     lc_trk_g2, lc_trk_g3, pgate, prog, purst, reset_b, s_r, vdd_cntl,
     wl );
output  carry_out;


input  cin2local, clk, clkb, prog, purst, s_r;

output [7:0]  slf_op;

inout [27:0]  bl;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;

input [15:0]  vdd_cntl;
input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  pgate;
input [7:0]  lc_trk_g1;
input [7:0]  lc_trk_g2;
input [7:0]  lc_trk_g3;
input [7:0]  lc_trk_g0;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;



lcmuxod3_0rev ILC_00 ( .clk(clk), .cbitb(cbitb[55:0]),
     .cbit(cbit[55:0]), .vdd_cntl(vdd_cntl[1:0]), .carry_in(cin),
     .op(slf_op[0]), .s_r(s_r), .purst(purst), .sp4_v_b({sp4_v_b[32],
     sp4_v_b[16], sp4_v_b[0]}), .reset_b(reset_b[1:0]),
     .sp4_h_r({sp4_h_r[32], sp4_h_r[16], sp4_h_r[0]}), .bl(bl[27:0]),
     .wl(wl[1:0]), .sp12_v_b({sp12_v_b[16], sp12_v_b[0]}),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], cin}),
     .sp4_r_v_b({sp4_r_v_b[33], sp4_r_v_b[17], sp4_r_v_b[1]}),
     .pgate(pgate[1:0]), .prog(prog), .sp12_h_r(sp12_h_r[8]),
     .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .carry_out(c_01));
lcmuxod3_0 ILC_03 ( .clk(clk), .vdd_cntl(vdd_cntl[7:6]),
     .carry_in(c_23), .op(slf_op[3]), .s_r(s_r), .purst(purst),
     .sp4_v_b({sp4_v_b[38], sp4_v_b[22], sp4_v_b[6]}),
     .reset_b(reset_b[7:6]), .sp4_h_r({sp4_h_r[38], sp4_h_r[22],
     sp4_h_r[6]}), .bl(bl[27:0]), .wl(wl[7:6]),
     .sp12_v_b({sp12_v_b[22], sp12_v_b[6]}), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], c_23}), .sp4_r_v_b({sp4_r_v_b[39],
     sp4_r_v_b[23], sp4_r_v_b[7]}), .pgate(pgate[7:6]), .prog(prog),
     .sp12_h_r(sp12_h_r[14]), .clkb(clkb), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .carry_out(c_34));
lcmuxod3_0 ILC_01 ( .clk(clk), .vdd_cntl(vdd_cntl[3:2]),
     .carry_in(c_01), .op(slf_op[1]), .s_r(s_r), .purst(purst),
     .sp4_v_b({sp4_v_b[34], sp4_v_b[18], sp4_v_b[2]}),
     .reset_b(reset_b[3:2]), .sp4_h_r({sp4_h_r[34], sp4_h_r[18],
     sp4_h_r[2]}), .bl(bl[27:0]), .wl(wl[3:2]),
     .sp12_v_b({sp12_v_b[18], sp12_v_b[2]}), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], c_01}), .sp4_r_v_b({sp4_r_v_b[35],
     sp4_r_v_b[19], sp4_r_v_b[3]}), .pgate(pgate[3:2]), .prog(prog),
     .sp12_h_r(sp12_h_r[10]), .clkb(clkb), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .carry_out(c_12));
lcmuxod3_0 ILC_02 ( .clk(clk), .vdd_cntl(vdd_cntl[5:4]),
     .carry_in(c_12), .op(slf_op[2]), .s_r(s_r), .purst(purst),
     .sp4_v_b({sp4_v_b[36], sp4_v_b[20], sp4_v_b[4]}),
     .reset_b(reset_b[5:4]), .sp4_h_r({sp4_h_r[36], sp4_h_r[20],
     sp4_h_r[4]}), .bl(bl[27:0]), .wl(wl[5:4]),
     .sp12_v_b({sp12_v_b[20], sp12_v_b[4]}), .min3({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], c_12}), .sp4_r_v_b({sp4_r_v_b[37],
     sp4_r_v_b[21], sp4_r_v_b[5]}), .pgate(pgate[5:4]), .prog(prog),
     .sp12_h_r(sp12_h_r[12]), .clkb(clkb), .min2({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .carry_out(c_23));
lcmuxod7_4 ILC_07 ( .clk(clk), .vdd_cntl(vdd_cntl[15:14]),
     .carry_in(c_67), .op(slf_op[7]), .s_r(s_r), .purst(purst),
     .sp4_v_b({sp4_v_b[46], sp4_v_b[30], sp4_v_b[14]}),
     .reset_b(reset_b[15:14]), .sp4_h_r({sp4_h_r[46], sp4_h_r[30],
     sp4_h_r[14]}), .bl(bl[27:0]), .wl(wl[15:14]),
     .sp12_v_b(sp12_v_b[14]), .sp12_h_r({sp12_h_r[22], sp12_h_r[6]}),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_67}),
     .carry_out(carry_out), .sp4_r_v_b({sp4_r_v_b[47], sp4_r_v_b[31],
     sp4_r_v_b[15]}), .pgate(pgate[15:14]), .prog(prog), .clkb(clkb),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}));
lcmuxod7_4 ILC_04 ( .clk(clk), .vdd_cntl(vdd_cntl[9:8]),
     .carry_in(c_34), .op(slf_op[4]), .s_r(s_r), .purst(purst),
     .sp4_v_b({sp4_v_b[40], sp4_v_b[24], sp4_v_b[8]}),
     .reset_b(reset_b[9:8]), .sp4_h_r({sp4_h_r[40], sp4_h_r[24],
     sp4_h_r[8]}), .bl(bl[27:0]), .wl(wl[9:8]), .sp12_v_b(sp12_v_b[8]),
     .sp12_h_r({sp12_h_r[16], sp12_h_r[0]}), .min3({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], c_34}), .carry_out(c_45),
     .sp4_r_v_b({sp4_r_v_b[41], sp4_r_v_b[25], sp4_r_v_b[9]}),
     .pgate(pgate[9:8]), .prog(prog), .clkb(clkb), .min2({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}));
lcmuxod7_4 ILC_05 ( .clk(clk), .vdd_cntl(vdd_cntl[11:10]),
     .carry_in(c_45), .op(slf_op[5]), .s_r(s_r), .purst(purst),
     .sp4_v_b({sp4_v_b[42], sp4_v_b[26], sp4_v_b[10]}),
     .reset_b(reset_b[11:10]), .sp4_h_r({sp4_h_r[42], sp4_h_r[26],
     sp4_h_r[10]}), .bl(bl[27:0]), .wl(wl[11:10]),
     .sp12_v_b(sp12_v_b[10]), .sp12_h_r({sp12_h_r[18], sp12_h_r[2]}),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_45}),
     .carry_out(c_56), .sp4_r_v_b({sp4_r_v_b[43], sp4_r_v_b[27],
     sp4_r_v_b[11]}), .pgate(pgate[11:10]), .prog(prog), .clkb(clkb),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}));
lcmuxod7_4 ILC_06 ( .clk(clk), .vdd_cntl(vdd_cntl[13:12]),
     .carry_in(c_56), .op(slf_op[6]), .s_r(s_r), .purst(purst),
     .sp4_v_b({sp4_v_b[44], sp4_v_b[28], sp4_v_b[12]}),
     .reset_b(reset_b[13:12]), .sp4_h_r({sp4_h_r[44], sp4_h_r[28],
     sp4_h_r[12]}), .bl(bl[27:0]), .wl(wl[13:12]),
     .sp12_v_b(sp12_v_b[12]), .sp12_h_r({sp12_h_r[20], sp12_h_r[4]}),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_56}),
     .carry_out(c_67), .sp4_r_v_b({sp4_r_v_b[45], sp4_r_v_b[29],
     sp4_r_v_b[13]}), .pgate(pgate[13:12]), .prog(prog), .clkb(clkb),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}));
mux_4carry Icarry_cnt ( .cin(cin2local), .lcl_cin(cin),
     .cbitb({cbitb[45], cbitb[48]}), .prog(prog), .cbit({cbit[45],
     cbit[48]}));

endmodule
// Library - leafcell, Cell - tielo, View - schematic
// LAST TIME SAVED: Jul  8 16:15:53 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module tielo ( tielo );
output  tielo;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M0 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));
nch_hvt  M1 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - leafcell, Cell - ltile4rev0, View - schematic
// LAST TIME SAVED: Jan 20 09:17:17 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module ltile4rev0 ( carry_out, cbit_colcntl, slf_op, bl, sp4_h_l,
     sp4_h_r, sp4_r_v_b, sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r,
     sp12_v_b, sp12_v_t, bnl_op, bnr_op, bot_op, carry_in, glb_netwk,
     lft_op, pgate, prog, purst, reset_b, rgt_op, tnl_op, tnr_op,
     top_op, vdd_cntl, wl );
output  carry_out;


input  carry_in, prog, purst;

output [7:0]  slf_op;
output [7:0]  cbit_colcntl;

inout [47:0]  sp4_v_t;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [23:0]  sp12_v_t;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_h_r;
inout [53:0]  bl;
inout [23:0]  sp12_v_b;

input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  glb_netwk;
input [7:0]  bot_op;
input [7:0]  top_op;
input [7:0]  bnl_op;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  wl;
input [15:0]  reset_b;
input [7:0]  bnr_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  lc_trk_g1;

wire  [7:0]  lc_trk_g3;

wire  [7:0]  lc_trk_g2;

wire  [1:0]  sp12_v_b_mid;

wire  [7:0]  lc_trk_g0;

wire  [3:0]  net_glb2local;

wire  [1:0]  sp12_h_r_mid;



gmux_sp12to4 Igmux_sp12to4 ( .reset_b({reset_b[14], reset_b[15],
     reset_b[12], reset_b[13], reset_b[10], reset_b[11], reset_b[8],
     reset_b[9], reset_b[6], reset_b[7], reset_b[4], reset_b[5],
     reset_b[2], reset_b[3], reset_b[0], reset_b[1]}),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .wl({wl[14], wl[15],
     wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4],
     wl[5], wl[2], wl[3], wl[0], wl[1]}), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .prog(progd), .lft_op(lft_op[7:0]),
     .bnr_op(bnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .lc_trk_g3(lc_trk_g3[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .bot_op(bot_op[7:0]), .glb2local(net_glb2local[3:0]),
     .sp12_v_b(sp12_v_b[23:0]), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[25:14]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]));
span4 Isp4_sw ( .pgate({pgate[14], pgate[15], pgate[12], pgate[13],
     pgate[10], pgate[11], pgate[8], pgate[9], pgate[6], pgate[7],
     pgate[4], pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .prog(progd), .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12],
     vdd_cntl[13], vdd_cntl[10], vdd_cntl[11], vdd_cntl[8],
     vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4], vdd_cntl[5],
     vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .reset_b({reset_b[14], reset_b[15], reset_b[12], reset_b[13],
     reset_b[10], reset_b[11], reset_b[8], reset_b[9], reset_b[6],
     reset_b[7], reset_b[4], reset_b[5], reset_b[2], reset_b[3],
     reset_b[0], reset_b[1]}), .wl({wl[14], wl[15], wl[12], wl[13],
     wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2],
     wl[3], wl[0], wl[1]}), .bl(bl[13:4]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_t(sp4_v_t[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp4_h_l(sp4_h_l[47:0]));
misc_module4rev0 I_misc ( .cbit_colcntl(cbit_colcntl[7:0]),
     .prog(progd), .lc_trk_g0(lc_trk_g0[5:0]),
     .glb_netwk(glb_netwk[7:0]), .lc_trk_g2(lc_trk_g2[5:0]),
     .lc_trk_g3(lc_trk_g3[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .S_R(s_r), .clkb(clkb), .bl(bl[3:0]), .clk(clk),
     .sp4(sp4_h_r[23:16]), .sp12({sp12_h_r[22], sp12_h_r[20],
     sp12_h_r[18], sp12_h_r[16], sp12_h_r[14], sp12_h_r[12],
     sp12_h_r[10], sp12_h_r[8]}), .reset_b({reset_b[14], reset_b[15],
     reset_b[12], reset_b[13], reset_b[10], reset_b[11], reset_b[8],
     reset_b[9], reset_b[6], reset_b[7], reset_b[4], reset_b[5],
     reset_b[2], reset_b[3], reset_b[0], reset_b[1]}),
     .b(sp12_v_b[1:0]), .r(sp12_h_r[1:0]), .m(sp12_v_b_mid[1:0]),
     .l(sp12_h_r_mid[1:0]), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12],
     vdd_cntl[13], vdd_cntl[10], vdd_cntl[11], vdd_cntl[8],
     vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4], vdd_cntl[5],
     vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .glb2local(net_glb2local[3:0]), .min2(glb_netwk[7:0]),
     .min1(glb_netwk[7:0]), .min0(glb_netwk[7:0]),
     .min3(glb_netwk[7:0]));
lccol_rev0 I_lccol_rev0 ( .s_r(s_r), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .reset_b({reset_b[14], reset_b[15], reset_b[12],
     reset_b[13], reset_b[10], reset_b[11], reset_b[8], reset_b[9],
     reset_b[6], reset_b[7], reset_b[4], reset_b[5], reset_b[2],
     reset_b[3], reset_b[0], reset_b[1]}), .prog(progd),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .purst(purst),
     .lc_trk_g3(lc_trk_g3[7:0]), .lc_trk_g2(lc_trk_g2[7:0]),
     .lc_trk_g1(lc_trk_g1[7:0]), .lc_trk_g0(lc_trk_g0[7:0]),
     .clkb(clkb), .clk(clk), .cin2local(carry_in),
     .slf_op(slf_op[7:0]), .carry_out(carry_out),
     .sp12_v_b(sp12_v_b[23:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .bl(bl[53:26]));
rm7  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
rm6  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm6  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm6  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm6  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm6  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm6  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm6  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm6  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm6  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm6  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm6  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm6  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm6  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm6  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm6  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm6  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm6  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm6  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm6  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm6  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm6  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm6  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm6  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm6  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
inv_hvt I89 ( .A(progb), .Y(progd));
inv_hvt I90 ( .A(prog), .Y(progb));

endmodule
// Library - leafcell, Cell - ice1f_array_LT_top, View - schematic
// LAST TIME SAVED: Jul  6 15:45:31 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module ice1f_array_LT_top ( carry_out, .glb_netwk_bo(glb_netwk_bot),
     .glb_netwk_to(glb_netwk_top), slf_op_01, slf_op_02, slf_op_03,
     slf_op_04, slf_op_05, slf_op_06, slf_op_07, slf_op_08, bl, pgate,
     reset_b, sp4_h_l_01, sp4_h_l_02, sp4_h_l_03, sp4_h_l_04,
     sp4_h_l_05, sp4_h_l_06, sp4_h_l_07, sp4_h_l_08, sp4_h_r_01,
     sp4_h_r_02, sp4_h_r_03, sp4_h_r_04, sp4_h_r_05, sp4_h_r_06,
     sp4_h_r_07, sp4_h_r_08, sp4_r_v_b_01, sp4_r_v_b_02, sp4_r_v_b_03,
     sp4_r_v_b_04, sp4_r_v_b_05, sp4_r_v_b_06, sp4_r_v_b_07,
     sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03, sp4_v_b_04,
     sp4_v_b_05, sp4_v_b_06, sp4_v_b_07, sp4_v_b_08, sp4_v_t_08,
     sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04, sp12_h_l_05,
     sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_r_01, sp12_h_r_02,
     sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06, sp12_h_r_07,
     sp12_h_r_08, sp12_v_b__01, sp12_v_t_08, vdd_cntl, wl, bnl_op_01,
     bnr_op_01, bot_op_01, carry_in, glb_netwk_col, lft_op_01,
     lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06, lft_op_07,
     lft_op_08, prog, purst, rgt_op_01, rgt_op_02, rgt_op_03,
     rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, tnl_op_08,
     tnr_op_08, top_op_08 );
output  carry_out;


input  carry_in, prog, purst;

output [7:0]  slf_op_08;
output [7:0]  slf_op_01;
output [7:0]  slf_op_02;
output [7:0]  slf_op_03;
output [7:0]  slf_op_06;
output [7:0]  glb_netwk_bot;
output [7:0]  glb_netwk_top;
output [7:0]  slf_op_04;
output [7:0]  slf_op_05;
output [7:0]  slf_op_07;

inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_h_r_06;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_r_v_b_04;
inout [47:0]  sp4_h_l_07;
inout [47:0]  sp4_h_l_08;
inout [47:0]  sp4_v_b_06;
inout [23:0]  sp12_h_l_06;
inout [47:0]  sp4_h_r_08;
inout [23:0]  sp12_h_l_03;
inout [23:0]  sp12_v_b__01;
inout [47:0]  sp4_h_l_06;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_h_r_04;
inout [47:0]  sp4_h_l_01;
inout [47:0]  sp4_v_b_03;
inout [23:0]  sp12_h_l_04;
inout [47:0]  sp4_r_v_b_02;
inout [47:0]  sp4_r_v_b_05;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_h_l_03;
inout [23:0]  sp12_h_r_06;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_v_b_07;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_v_b_02;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_v_b_05;
inout [23:0]  sp12_h_l_05;
inout [127:0]  vdd_cntl;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_h_l_04;
inout [23:0]  sp12_h_l_08;
inout [127:0]  wl;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_v_b_01;
inout [23:0]  sp12_h_r_04;
inout [23:0]  sp12_v_t_08;
inout [47:0]  sp4_h_l_02;
inout [23:0]  sp12_h_r_05;
inout [23:0]  sp12_h_r_08;
inout [53:0]  bl;
inout [47:0]  sp4_h_l_05;
inout [127:0]  reset_b;
inout [47:0]  sp4_h_r_02;
inout [127:0]  pgate;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_v_t_08;
inout [23:0]  sp12_h_l_07;

input [7:0]  bnr_op_01;
input [7:0]  rgt_op_06;
input [7:0]  rgt_op_05;
input [7:0]  lft_op_08;
input [7:0]  bnl_op_01;
input [7:0]  lft_op_03;
input [7:0]  lft_op_01;
input [7:0]  tnr_op_08;
input [7:0]  rgt_op_01;
input [7:0]  rgt_op_02;
input [7:0]  bot_op_01;
input [7:0]  rgt_op_04;
input [7:0]  lft_op_04;
input [7:0]  rgt_op_08;
input [7:0]  glb_netwk_col;
input [7:0]  lft_op_07;
input [7:0]  lft_op_05;
input [7:0]  lft_op_02;
input [7:0]  top_op_08;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_03;
input [7:0]  tnl_op_08;
input [7:0]  lft_op_06;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net572;

wire  [0:7]  net336;

wire  [0:23]  net346;

wire  [7:0]  colbuf_cntl_b;

wire  [7:0]  colbuf_cntl_t;

wire  [0:23]  net491;

wire  [0:23]  net375;

wire  [0:7]  net365;

wire  [0:7]  net577;

wire  [0:23]  net462;

wire  [0:7]  net575;

wire  [0:23]  net433;

wire  [0:23]  net404;

wire  [0:23]  net549;

wire  [0:7]  net571;



clk_colbuf1kx8 I_clk_colbuf1kx8_t ( .colbuf_cntl(colbuf_cntl_t[7:0]),
     .col_clk(glb_netwk_top[7:0]), .clk_in(glb_netwk_col[7:0]));
clk_colbuf1kx8 I_clk_colbuf12kx8_b ( .colbuf_cntl(colbuf_cntl_b[7:0]),
     .col_clk(glb_netwk_bot[7:0]), .clk_in(glb_netwk_col[7:0]));
ltile4rev0 I_LT06 ( .cbit_colcntl(net336[0:7]), .prog(prog),
     .carry_out(net338), .lft_op(lft_op_06[7:0]),
     .sp12_h_l(sp12_h_l_06[23:0]), .sp4_h_l(sp4_h_l_06[47:0]),
     .sp4_v_b(sp4_v_b_06[47:0]), .sp12_v_b(net433[0:23]),
     .sp12_h_r(sp12_h_r_06[23:0]), .sp4_h_r(sp4_h_r_06[47:0]),
     .sp12_v_t(net346[0:23]), .sp4_v_t(sp4_v_b_07[47:0]),
     .sp4_r_v_b(sp4_r_v_b_06[47:0]), .wl(wl[95:80]),
     .top_op(slf_op_07[7:0]), .rgt_op(rgt_op_06[7:0]),
     .bot_op(slf_op_05[7:0]), .bl(bl[53:0]), .reset_b(reset_b[95:80]),
     .vdd_cntl(vdd_cntl[95:80]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net425), .purst(purst), .slf_op(slf_op_06[7:0]),
     .pgate(pgate[95:80]), .bnr_op(rgt_op_05[7:0]),
     .bnl_op(lft_op_05[7:0]), .tnr_op(rgt_op_07[7:0]),
     .tnl_op(lft_op_07[7:0]));
ltile4rev0 I_LT03 ( .cbit_colcntl(net365[0:7]), .prog(prog),
     .carry_out(net367), .lft_op(lft_op_03[7:0]),
     .sp12_h_l(sp12_h_l_03[23:0]), .sp4_h_l(sp4_h_l_03[47:0]),
     .sp4_v_b(sp4_v_b_03[47:0]), .sp12_v_b(net491[0:23]),
     .sp12_h_r(sp12_h_r_03[23:0]), .sp4_h_r(sp4_h_r_03[47:0]),
     .sp12_v_t(net375[0:23]), .sp4_v_t(sp4_v_b_04[47:0]),
     .sp4_r_v_b(sp4_r_v_b_03[47:0]), .wl(wl[47:32]),
     .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net483), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4rev0 I_LT04 ( .cbit_colcntl(colbuf_cntl_b[7:0]), .prog(prog),
     .carry_out(net396), .lft_op(lft_op_04[7:0]),
     .sp12_h_l(sp12_h_l_04[23:0]), .sp4_h_l(sp4_h_l_04[47:0]),
     .sp4_v_b(sp4_v_b_04[47:0]), .sp12_v_b(net375[0:23]),
     .sp12_h_r(sp12_h_r_04[23:0]), .sp4_h_r(sp4_h_r_04[47:0]),
     .sp12_v_t(net404[0:23]), .sp4_v_t(sp4_v_b_05[47:0]),
     .sp4_r_v_b(sp4_r_v_b_04[47:0]), .wl(wl[63:48]),
     .top_op(slf_op_05[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net367), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(rgt_op_05[7:0]),
     .tnl_op(lft_op_05[7:0]));
ltile4rev0 I_LT05 ( .cbit_colcntl(colbuf_cntl_t[7:0]), .prog(prog),
     .carry_out(net425), .lft_op(lft_op_05[7:0]),
     .sp12_h_l(sp12_h_l_05[23:0]), .sp4_h_l(sp4_h_l_05[47:0]),
     .sp4_v_b(sp4_v_b_05[47:0]), .sp12_v_b(net404[0:23]),
     .sp12_h_r(sp12_h_r_05[23:0]), .sp4_h_r(sp4_h_r_05[47:0]),
     .sp12_v_t(net433[0:23]), .sp4_v_t(sp4_v_b_06[47:0]),
     .sp4_r_v_b(sp4_r_v_b_05[47:0]), .wl(wl[79:64]),
     .top_op(slf_op_06[7:0]), .rgt_op(rgt_op_05[7:0]),
     .bot_op(slf_op_04[7:0]), .bl(bl[53:0]), .reset_b(reset_b[79:64]),
     .vdd_cntl(vdd_cntl[79:64]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net396), .purst(purst), .slf_op(slf_op_05[7:0]),
     .pgate(pgate[79:64]), .bnr_op(rgt_op_04[7:0]),
     .bnl_op(lft_op_04[7:0]), .tnr_op(rgt_op_06[7:0]),
     .tnl_op(lft_op_06[7:0]));
ltile4rev0 I_LT01 ( .cbit_colcntl(net577[0:7]), .prog(prog),
     .carry_out(net454), .lft_op(lft_op_01[7:0]),
     .sp12_h_l(sp12_h_l_01[23:0]), .sp4_h_l(sp4_h_l_01[47:0]),
     .sp4_v_b(sp4_v_b_01[47:0]), .sp12_v_b(sp12_v_b__01[23:0]),
     .sp12_h_r(sp12_h_r_01[23:0]), .sp4_h_r(sp4_h_r_01[47:0]),
     .sp12_v_t(net462[0:23]), .sp4_v_t(sp4_v_b_02[47:0]),
     .sp4_r_v_b(sp4_r_v_b_01[47:0]), .wl(wl[15:0]),
     .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4rev0 I_LT02 ( .cbit_colcntl(net572[0:7]), .prog(prog),
     .carry_out(net483), .lft_op(lft_op_02[7:0]),
     .sp12_h_l(sp12_h_l_02[23:0]), .sp4_h_l(sp4_h_l_02[47:0]),
     .sp4_v_b(sp4_v_b_02[47:0]), .sp12_v_b(net462[0:23]),
     .sp12_h_r(sp12_h_r_02[23:0]), .sp4_h_r(sp4_h_r_02[47:0]),
     .sp12_v_t(net491[0:23]), .sp4_v_t(sp4_v_b_03[47:0]),
     .sp4_r_v_b(sp4_r_v_b_02[47:0]), .wl(wl[31:16]),
     .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net454), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));
ltile4rev0 I_LT08 ( .cbit_colcntl(net575[0:7]), .prog(prog),
     .carry_out(carry_out), .lft_op(lft_op_08[7:0]),
     .sp12_h_l(sp12_h_l_08[23:0]), .sp4_h_l(sp4_h_l_08[47:0]),
     .sp4_v_b(sp4_v_b_08[47:0]), .sp12_v_b(net549[0:23]),
     .sp12_h_r(sp12_h_r_08[23:0]), .sp4_h_r(sp4_h_r_08[47:0]),
     .sp12_v_t(sp12_v_t_08[23:0]), .sp4_v_t(sp4_v_t_08[47:0]),
     .sp4_r_v_b(sp4_r_v_b_08[47:0]), .wl(wl[127:112]),
     .top_op(top_op_08[7:0]), .rgt_op(rgt_op_08[7:0]),
     .bot_op(slf_op_07[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[127:112]), .vdd_cntl(vdd_cntl[127:112]),
     .glb_netwk(glb_netwk_top[7:0]), .carry_in(net541), .purst(purst),
     .slf_op(slf_op_08[7:0]), .pgate(pgate[127:112]),
     .bnr_op(rgt_op_07[7:0]), .bnl_op(lft_op_07[7:0]),
     .tnr_op(tnr_op_08[7:0]), .tnl_op(tnl_op_08[7:0]));
ltile4rev0 I_LT07 ( .cbit_colcntl(net571[0:7]), .prog(prog),
     .carry_out(net541), .lft_op(lft_op_07[7:0]),
     .sp12_h_l(sp12_h_l_07[23:0]), .sp4_h_l(sp4_h_l_07[47:0]),
     .sp4_v_b(sp4_v_b_07[47:0]), .sp12_v_b(net346[0:23]),
     .sp12_h_r(sp12_h_r_07[23:0]), .sp4_h_r(sp4_h_r_07[47:0]),
     .sp12_v_t(net549[0:23]), .sp4_v_t(sp4_v_b_08[47:0]),
     .sp4_r_v_b(sp4_r_v_b_07[47:0]), .wl(wl[111:96]),
     .top_op(slf_op_08[7:0]), .rgt_op(rgt_op_07[7:0]),
     .bot_op(slf_op_06[7:0]), .bl(bl[53:0]), .reset_b(reset_b[111:96]),
     .vdd_cntl(vdd_cntl[111:96]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net338), .purst(purst), .slf_op(slf_op_07[7:0]),
     .pgate(pgate[111:96]), .bnr_op(rgt_op_06[7:0]),
     .bnl_op(lft_op_06[7:0]), .tnr_op(rgt_op_08[7:0]),
     .tnl_op(lft_op_08[7:0]));

endmodule
// Library - leafcell, Cell - bram_routing_tracks4rev12, View -
//schematic
// LAST TIME SAVED: Jan 29 16:25:42 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_routing_tracks4rev12 ( cbit_colcntl, clk, lc_trk_g0,
     lc_trk_g1, lc_trk_g2, lc_trk_g3, s_r, bl, sp4_h_l, sp4_h_r,
     sp4_r_v_b, sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r, sp12_v_b,
     sp12_v_t, bnl_op, bnr_op, bot_op, glb_netwk, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );
output  clk, s_r;


input  prog;

output [7:0]  cbit_colcntl;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g3;
output [7:0]  lc_trk_g1;

inout [47:0]  sp4_v_t;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_l;
inout [25:0]  bl;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_v_t;

input [7:0]  bnl_op;
input [7:0]  glb_netwk;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  slf_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
input [15:0]  reset_b;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [15:0]  vdd_cntl;
input [7:0]  top_op;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net_glb2local;

wire  [1:0]  sp12_h_r_mid;

wire  [1:0]  sp12_v_b_mid;



gmux_sp12to4 Igmux_sp12to4 ( .reset_b(reset_b[15:0]),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .wl(wl[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .prog(progd), .lft_op(lft_op[7:0]),
     .bnr_op(bnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .lc_trk_g3(lc_trk_g3[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .bot_op(bot_op[7:0]), .glb2local(net_glb2local[3:0]),
     .sp12_v_b(sp12_v_b[23:0]), .pgate(pgate[15:0]), .bl(bl[25:14]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_r(sp4_h_r[47:0]));
span4 Isp4_sw ( .pgate(pgate[15:0]), .prog(progd),
     .vdd_cntl(vdd_cntl[15:0]), .reset_b(reset_b[15:0]), .wl(wl[15:0]),
     .bl(bl[13:4]), .sp4_h_r(sp4_h_r[47:0]), .sp4_v_t(sp4_v_t[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_l(sp4_h_l[47:0]));
misc_module4rev0 I_misc ( .cbit_colcntl(cbit_colcntl[7:0]),
     .prog(progd), .lc_trk_g0(lc_trk_g0[5:0]),
     .glb_netwk(glb_netwk[7:0]), .lc_trk_g2(lc_trk_g2[5:0]),
     .lc_trk_g3(lc_trk_g3[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .wl(wl[15:0]), .S_R(s_r), .clkb(net147), .bl(bl[3:0]), .clk(clk),
     .sp4(sp4_h_r[23:16]), .sp12({sp12_h_r[22], sp12_h_r[20],
     sp12_h_r[18], sp12_h_r[16], sp12_h_r[14], sp12_h_r[12],
     sp12_h_r[10], sp12_h_r[8]}), .reset_b(reset_b[15:0]),
     .b(sp12_v_b[1:0]), .r(sp12_h_r[1:0]), .m(sp12_v_b_mid[1:0]),
     .l(sp12_h_r_mid[1:0]), .pgate(pgate[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb2local(net_glb2local[3:0]),
     .min2(glb_netwk[7:0]), .min1(glb_netwk[7:0]),
     .min0(glb_netwk[7:0]), .min3(glb_netwk[7:0]));
rm7  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
rm6  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm6  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm6  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm6  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm6  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm6  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm6  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm6  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm6  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm6  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm6  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm6  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm6  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm6  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm6  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm6  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm6  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm6  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm6  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm6  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm6  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm6  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm6  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm6  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
inv_hvt I89 ( .A(progb), .Y(progd));
inv_hvt I90 ( .A(prog), .Y(progb));

endmodule
// Library - leafcell, Cell - bram_bufferx6, View - schematic
// LAST TIME SAVED: Jun 25 13:45:32 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_bufferx6 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jun  5 11:34:46 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module leafcell_ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - leafcell, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:59 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module ml_mux2_hvt_schematic ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - leafcell, Cell - bram_dff_mux, View - schematic
// LAST TIME SAVED: Jul 25 16:06:22 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_dff_mux ( q, bm_q, bm_sdi, ce, clk, rcapmux_en, rst );
output  q;

input  bm_q, bm_sdi, ce, clk, rcapmux_en, rst;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



leafcell_ml_dff_schematic I2 ( .R(rst), .D(net020), .CLK(clk),
     .QN(net10), .Q(q));
ml_mux2_hvt_schematic I5 ( .in1(net14), .in0(q), .out(net020),
     .sel(ce));
ml_mux2_hvt_schematic I1 ( .in1(bm_q), .in0(bm_sdi), .out(net14),
     .sel(rcapmux_en));

endmodule
// Library - leafcell, Cell - bram_4k_sr, View - schematic
// LAST TIME SAVED: Aug 15 17:41:16 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4k_sr ( bm_dm, bm_sweb, clk, rcapmux_en, rst, bm_q, bm_sdi,
     wdummymux_en );

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[0]), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));

endmodule
// Library - leafcell, Cell - rf_4k, View - schematic
// LAST TIME SAVED: Aug 15 17:39:16 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module rf_4k ( Q, AA, AB, AMA, AMB, BIST, BWEB, BWEBM, CLKR, CLKW, D,
     DM, REB, REBM, WEB, WEBM );

input  BIST, CLKR, CLKW, REB, REBM, WEB, WEBM;

output [15:0]  Q;

input [7:0]  AMA;
input [15:0]  BWEBM;
input [15:0]  DM;
input [7:0]  AA;
input [15:0]  D;
input [15:0]  BWEB;
input [7:0]  AMB;
input [7:0]  AB;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - leafcell, Cell - bram_4k, View - schematic
// LAST TIME SAVED: Aug 15 17:44:47 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4k ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr, bm_clkw,
     bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk, bm_sclkrw,
     bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_sa;
input [7:0]  bm_ab;
input [7:0]  bm_aa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [14:0]  bm_dm;



tielo I15 ( .tielo(net101));
tielo I18 ( .tielo(net102));
bram_4k_sr I12 ( .bm_dm({bm_sdo, bm_dm[14:0]}), .rst(net102),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM({bm_sdo, bm_dm[14:0]}), .WEBM(bm_sweb), .WEB(web),
     .REBM(bm_sreb), .REB(reb), .D(bm_d[15:0]), .CLKW(net81),
     .CLKR(net79), .BWEBM({net101, net101, net101, net101, net101,
     net101, net101, net101, net101, net101, net101, net101, net101,
     net101, net101, net101}), .BWEB(bm_bweb[15:0]), .BIST(bm_init),
     .AMB(bm_sa[7:0]), .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]),
     .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net97), .out(net79));
bram_bufferx6 I8 ( .in(net93), .out(net81));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net93), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net97), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - misc, Cell - ml_mux3_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:41 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_mux3_hvt ( out, in0, in1, in2, sel );
output  out;

input  in0, in1, in2;

input [3:0]  sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I25 ( .A(sel[2]), .Y(net26));
inv_hvt I24 ( .A(sel[1]), .Y(net28));
inv_hvt I21 ( .A(sel[0]), .Y(net30));
txgate_hvt I23 ( .in(in1), .out(out), .pp(net28), .nn(sel[1]));
txgate_hvt I20 ( .in(in0), .out(out), .pp(net30), .nn(sel[0]));
txgate_hvt I26 ( .in(in2), .out(out), .pp(net26), .nn(sel[2]));
nch_hvt  MN19 ( .D(out), .B(gnd_), .G(sel[3]), .S(gnd_));

endmodule
// Library - leafcell, Cell - bram_bufferx1, View - schematic
// LAST TIME SAVED: Jun 14 08:59:24 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_bufferx1 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I0 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(in), .Y(net6));

endmodule
// Library - leafcell, Cell - bram_4k_buffer, View - schematic
// LAST TIME SAVED: Oct  6 13:53:19 2008
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4k_buffer ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;

input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



tielo I22 ( .tielo(net055));
bram_bufferx1 I15 ( .in(net055), .out(net49));
bram_bufferx1 I16 ( .in(net49), .out(net52));
bram_bufferx1 I17 ( .in(net52), .out(net53));
bram_bufferx1 I18 ( .in(net53), .out(net55));
bram_bufferx6 I14 ( .in(bm_sdo_i), .out(bm_sdo_o));
bram_bufferx6 I6 ( .in(bm_sdi_i), .out(bm_sdi_o));
bram_bufferx6 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx6 I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx6 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx6 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx6 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx6 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx6 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx6 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx6 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx6 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx6 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx6 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx6 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx6 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx6 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - bram_4kbank_pbuffer_bot, View - schematic
// LAST TIME SAVED: Aug 24 17:32:39 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4kbank_pbuffer_bot ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sclkrw_o;
output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;

input [15:0]  bm_d;
input [15:0]  bm_bweb;
input [1:0]  bm_sweb_i;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sdo_i;
input [7:0]  bm_ab;
input [1:0]  bm_sclkrw_i;
input [7:0]  bm_sa_i;
input [7:0]  bm_aa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o[0]), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i[0]), .bm_sclkrw_o(bm_sclkrw_o[0]),
     .bm_sdi_o(bm_sdi_o[0]), .bm_sdi_i(bm_sdi_i[0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));

endmodule
// Library - leafcell, Cell - bram_4k_inmux3_0, View - schematic
// LAST TIME SAVED: Aug 23 11:45:13 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4k_inmux3_0 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_h_r;

input  op, prog;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_v_b;

input [15:0]  min3;
input [15:0]  min0;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [15:0]  min1;
input [15:0]  bl;
input [15:0]  min2;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [31:0]  cbitb;

wire  [31:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
odrv12_30 Iodrv74 ( .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
in_mux in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12], cbit[13],
     cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux7_4, View - schematic
// LAST TIME SAVED: Aug 23 11:44:11 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4k_inmux7_4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_v_b;

input  op, prog;

output [1:0]  sp12_h_r;
output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;

input [15:0]  min3;
input [15:0]  min0;
input [15:0]  bl;
input [1:0]  vdd_cntl;
input [15:0]  min1;
input [1:0]  wl;
input [1:0]  pgate;
input [15:0]  min2;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [31:0]  cbit;

wire  [31:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
odrv12_74 Iodrv74 ( .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .sp12_v_b(sp12_v_b),
     .sp12_h_r(sp12_h_r[1:0]));
in_mux in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12], cbit[13],
     cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux_8x4, View - schematic
// LAST TIME SAVED: Aug 29 16:20:56 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4k_inmux_8x4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, op, pgate, prog, reset_b, vdd_cntl, wl );

input  prog;

output [23:0]  sp4_r_v_b;
output [23:0]  sp4_h_r;
output [7:0]  in3;
output [7:0]  in2;
output [7:0]  in1;
output [11:0]  sp12_v_b;
output [11:0]  sp12_h_r;
output [23:0]  sp4_v_b;
output [7:0]  in0;

input [15:0]  bl;
input [7:0]  op;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g2;
input [15:0]  reset_b;
input [7:0]  lc_trk_g1;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [7:0]  lc_trk_g3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_4k_inmux3_0 I3 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[3]), .sp12_v_b(sp12_v_b[7:6]), .wl(wl[7:6]),
     .reset_b(reset_b[7:6]), .prog(progd), .pgate(pgate[7:6]),
     .op(op[3]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[11:9]), .sp4_r_v_b(sp4_r_v_b[11:9]),
     .sp4_h_r(sp4_h_r[11:9]), .in3(in3[3]), .in2(in2[3]), .in1(in1[3]),
     .in0(in0[3]));
bram_4k_inmux3_0 I2 ( .vdd_cntl(vdd_cntl[5:4]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[2]), .sp12_v_b(sp12_v_b[5:4]), .wl(wl[5:4]),
     .reset_b(reset_b[5:4]), .prog(progd), .pgate(pgate[5:4]),
     .op(op[2]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[8:6]), .sp4_r_v_b(sp4_r_v_b[8:6]),
     .sp4_h_r(sp4_h_r[8:6]), .in3(in3[2]), .in2(in2[2]), .in1(in1[2]),
     .in0(in0[2]));
bram_4k_inmux3_0 I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[1]), .sp12_v_b(sp12_v_b[3:2]), .wl(wl[3:2]),
     .reset_b(reset_b[3:2]), .prog(progd), .pgate(pgate[3:2]),
     .op(op[1]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[5:3]), .sp4_r_v_b(sp4_r_v_b[5:3]),
     .sp4_h_r(sp4_h_r[5:3]), .in3(in3[1]), .in2(in2[1]), .in1(in1[1]),
     .in0(in0[1]));
bram_4k_inmux3_0 I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[0]), .sp12_v_b(sp12_v_b[1:0]), .wl(wl[1:0]),
     .reset_b(reset_b[1:0]), .prog(progd), .pgate(pgate[1:0]),
     .op(op[0]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_r_v_b(sp4_r_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .in3(in3[0]), .in2(in2[0]), .in1(in1[0]),
     .in0(in0[0]));
tiehi I10 ( .tiehi(tiehi));
bram_4k_inmux7_4 I6 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[15:0]),
     .wl(wl[13:12]), .reset_b(reset_b[13:12]), .prog(progd),
     .pgate(pgate[13:12]), .op(op[6]), .min3({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp12_v_b(sp12_v_b[10]), .sp12_h_r(sp12_h_r[9:8]),
     .sp4_v_b(sp4_v_b[20:18]), .sp4_r_v_b(sp4_r_v_b[20:18]),
     .sp4_h_r(sp4_h_r[20:18]), .in3(in3[6]), .in2(in2[6]),
     .in1(in1[6]), .in0(in0[6]));
bram_4k_inmux7_4 I5 ( .vdd_cntl(vdd_cntl[11:10]), .bl(bl[15:0]),
     .wl(wl[11:10]), .reset_b(reset_b[11:10]), .prog(progd),
     .pgate(pgate[11:10]), .op(op[5]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[9]), .sp12_h_r(sp12_h_r[7:6]),
     .sp4_v_b(sp4_v_b[17:15]), .sp4_r_v_b(sp4_r_v_b[17:15]),
     .sp4_h_r(sp4_h_r[17:15]), .in3(in3[5]), .in2(in2[5]),
     .in1(in1[5]), .in0(in0[5]));
bram_4k_inmux7_4 I4 ( .vdd_cntl(vdd_cntl[9:8]), .bl(bl[15:0]),
     .wl(wl[9:8]), .reset_b(reset_b[9:8]), .prog(progd),
     .pgate(pgate[9:8]), .op(op[4]), .min3({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .sp12_v_b(sp12_v_b[8]),
     .sp12_h_r(sp12_h_r[5:4]), .sp4_v_b(sp4_v_b[14:12]),
     .sp4_r_v_b(sp4_r_v_b[14:12]), .sp4_h_r(sp4_h_r[14:12]),
     .in3(in3[4]), .in2(in2[4]), .in1(in1[4]), .in0(in0[4]));
bram_4k_inmux7_4 I7 ( .vdd_cntl(vdd_cntl[15:14]), .bl(bl[15:0]),
     .wl(wl[15:14]), .reset_b(reset_b[15:14]), .prog(progd),
     .pgate(pgate[15:14]), .op(op[7]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[11]), .sp12_h_r(sp12_h_r[11:10]),
     .sp4_v_b(sp4_v_b[23:21]), .sp4_r_v_b(sp4_r_v_b[23:21]),
     .sp4_h_r(sp4_h_r[23:21]), .in3(in3[7]), .in2(in2[7]),
     .in1(in1[7]), .in0(in0[7]));
inv_hvt I81 ( .A(prog), .Y(progb));
inv_hvt I82 ( .A(progb), .Y(progd));

endmodule
// Library - leafcell, Cell - bram_4kprouting_bbank, View - schematic
// LAST TIME SAVED: Jan  8 09:21:37 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4kprouting_bbank ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, cbit_colcntl, slf_op_bot, slf_op_top, bl,
     sp4_h_l_bot, sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [7:0]  cbit_colcntl;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sclkrw_o;

inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_h_l_bot;
inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_h_l_top;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_r_v_b_top;
inout [41:0]  bl;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_r_v_b_bot;

input [7:0]  bm_sa_i;
input [7:0]  tnr_op_bot;
input [1:0]  bm_sweb_i;
input [7:0]  bnl_op_bot;
input [7:0]  glb_netwk;
input [7:0]  tnl_op_top;
input [7:0]  rgt_op_top;
input [15:0]  reset_b_bot;
input [1:0]  bm_sclkrw_i;
input [7:0]  bnr_op_bot;
input [7:0]  top_op_top;
input [7:0]  bnl_op_top;
input [7:0]  rgt_op_bot;
input [7:0]  bnr_op_top;
input [15:0]  pgate_bot;
input [1:0]  bm_sdi_i;
input [7:0]  lft_op_top;
input [15:0]  pgate_top;
input [15:0]  wl_bot;
input [15:0]  vdd_cntl_top;
input [15:0]  reset_b_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  bot_op_bot;
input [7:0]  tnr_op_top;
input [1:0]  bm_sdo_i;
input [7:0]  tnl_op_bot;
input [7:0]  lft_op_bot;
input [15:0]  wl_top;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net226;

wire  [0:7]  net261;

wire  [0:7]  net229;

wire  [0:7]  net343;

wire  [0:7]  net227;

wire  [0:7]  net259;

wire  [15:0]  bm_bweb;

wire  [0:7]  net228;

wire  [0:7]  net260;

wire  [7:0]  in2_bot;

wire  [0:7]  net322;

wire  [0:7]  net258;

wire  [0:7]  net0239;

wire  [23:0]  sp12_v_b_top;

wire  [15:0]  bm_d;

wire  [7:0]  in2_top;



bram_routing_tracks4rev12 I_bot ( .cbit_colcntl(cbit_colcntl[7:0]),
     .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15], vdd_cntl_bot[12],
     vdd_cntl_bot[13], vdd_cntl_bot[10], vdd_cntl_bot[11],
     vdd_cntl_bot[8], vdd_cntl_bot[9], vdd_cntl_bot[6],
     vdd_cntl_bot[7], vdd_cntl_bot[4], vdd_cntl_bot[5],
     vdd_cntl_bot[2], vdd_cntl_bot[3], vdd_cntl_bot[0],
     vdd_cntl_bot[1]}), .s_r(net210), .wl({wl_bot[14], wl_bot[15],
     wl_bot[12], wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8],
     wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2],
     wl_bot[3], wl_bot[0], wl_bot[1]}), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net226[0:7]),
     .lc_trk_g2(net227[0:7]), .lc_trk_g1(net228[0:7]),
     .lc_trk_g0(net229[0:7]), .clk(net230),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev12 I_top ( .cbit_colcntl(net0239[0:7]),
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .s_r(net242), .wl({wl_top[14], wl_top[15],
     wl_top[12], wl_top[13], wl_top[10], wl_top[11], wl_top[8],
     wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2],
     wl_top[3], wl_top[0], wl_top[1]}), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net258[0:7]),
     .lc_trk_g2(net259[0:7]), .lc_trk_g1(net260[0:7]),
     .lc_trk_g0(net261[0:7]), .clk(net262),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbank_pbuffer_bot I_bram_4kbank_pbuffer_bot (
     .bm_q({slf_op_top[7:0], slf_op_bot[7:0]}),
     .bm_sdo_i(bm_sdo_i[1:0]), .bm_sdi_o(bm_sdi_o[1:0]),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sdi_i(bm_sdi_i[1:0]),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .bm_sweb_i(bm_sweb_i[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sweb_o(bm_sweb_o[1:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_init_i(bm_init_i),
     .bm_ren(net242), .bm_wen(net210), .bm_d(bm_d[15:0]),
     .bm_clkr(net262), .bm_clkw(net230), .bm_bweb(bm_bweb[15:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_ab(net343[0:7]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sreb_i(bm_sreb_i), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_aa(net322[0:7]), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I_inmux_8x4_b ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}),
     .bl(bl[41:26]), .wl({wl_bot[14], wl_bot[15], wl_bot[12],
     wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8], wl_bot[9],
     wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2], wl_bot[3],
     wl_bot[0], wl_bot[1]}), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .op(slf_op_bot[7:0]), .lc_trk_g3(net226[0:7]),
     .lc_trk_g2(net227[0:7]), .lc_trk_g1(net228[0:7]),
     .lc_trk_g0(net229[0:7]), .sp12_h_r({sp12_h_r_bot[22],
     sp12_h_r_bot[6], sp12_h_r_bot[20], sp12_h_r_bot[4],
     sp12_h_r_bot[18], sp12_h_r_bot[2], sp12_h_r_bot[16],
     sp12_h_r_bot[0], sp12_h_r_bot[14], sp12_h_r_bot[12],
     sp12_h_r_bot[10], sp12_h_r_bot[8]}), .sp4_v_b({sp4_v_b_bot[46],
     sp4_v_b_bot[30], sp4_v_b_bot[14], sp4_v_b_bot[44],
     sp4_v_b_bot[28], sp4_v_b_bot[12], sp4_v_b_bot[42],
     sp4_v_b_bot[26], sp4_v_b_bot[10], sp4_v_b_bot[40],
     sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38], sp4_v_b_bot[22],
     sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20], sp4_v_b_bot[4],
     sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2], sp4_v_b_bot[32],
     sp4_v_b_bot[16], sp4_v_b_bot[0]}), .sp4_r_v_b({sp4_r_v_b_bot[47],
     sp4_r_v_b_bot[31], sp4_r_v_b_bot[15], sp4_r_v_b_bot[45],
     sp4_r_v_b_bot[29], sp4_r_v_b_bot[13], sp4_r_v_b_bot[43],
     sp4_r_v_b_bot[27], sp4_r_v_b_bot[11], sp4_r_v_b_bot[41],
     sp4_r_v_b_bot[25], sp4_r_v_b_bot[9], sp4_r_v_b_bot[39],
     sp4_r_v_b_bot[23], sp4_r_v_b_bot[7], sp4_r_v_b_bot[37],
     sp4_r_v_b_bot[21], sp4_r_v_b_bot[5], sp4_r_v_b_bot[35],
     sp4_r_v_b_bot[19], sp4_r_v_b_bot[3], sp4_r_v_b_bot[33],
     sp4_r_v_b_bot[17], sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46],
     sp4_h_r_bot[30], sp4_h_r_bot[14], sp4_h_r_bot[44],
     sp4_h_r_bot[28], sp4_h_r_bot[12], sp4_h_r_bot[42],
     sp4_h_r_bot[26], sp4_h_r_bot[10], sp4_h_r_bot[40],
     sp4_h_r_bot[24], sp4_h_r_bot[8], sp4_h_r_bot[38], sp4_h_r_bot[22],
     sp4_h_r_bot[6], sp4_h_r_bot[36], sp4_h_r_bot[20], sp4_h_r_bot[4],
     sp4_h_r_bot[34], sp4_h_r_bot[18], sp4_h_r_bot[2], sp4_h_r_bot[32],
     sp4_h_r_bot[16], sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]),
     .in2(in2_bot[7:0]), .in1(bm_d[7:0]), .in0(net322[0:7]),
     .sp12_v_b({sp12_v_b_bot[14], sp12_v_b_bot[12], sp12_v_b_bot[10],
     sp12_v_b_bot[8], sp12_v_b_bot[22], sp12_v_b_bot[6],
     sp12_v_b_bot[20], sp12_v_b_bot[4], sp12_v_b_bot[18],
     sp12_v_b_bot[2], sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I_inmux_8x4_t ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}),
     .bl(bl[41:26]), .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12],
     sp12_v_b_top[10], sp12_v_b_top[8], sp12_v_b_top[22],
     sp12_v_b_top[6], sp12_v_b_top[20], sp12_v_b_top[4],
     sp12_v_b_top[18], sp12_v_b_top[2], sp12_v_b_top[16],
     sp12_v_b_top[0]}), .wl({wl_top[14], wl_top[15], wl_top[12],
     wl_top[13], wl_top[10], wl_top[11], wl_top[8], wl_top[9],
     wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2], wl_top[3],
     wl_top[0], wl_top[1]}), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .op(slf_op_top[7:0]), .lc_trk_g3(net258[0:7]),
     .lc_trk_g2(net259[0:7]), .lc_trk_g1(net260[0:7]),
     .lc_trk_g0(net261[0:7]), .sp12_h_r({sp12_h_r_top[22],
     sp12_h_r_top[6], sp12_h_r_top[20], sp12_h_r_top[4],
     sp12_h_r_top[18], sp12_h_r_top[2], sp12_h_r_top[16],
     sp12_h_r_top[0], sp12_h_r_top[14], sp12_h_r_top[12],
     sp12_h_r_top[10], sp12_h_r_top[8]}), .sp4_v_b({sp4_v_b_top[46],
     sp4_v_b_top[30], sp4_v_b_top[14], sp4_v_b_top[44],
     sp4_v_b_top[28], sp4_v_b_top[12], sp4_v_b_top[42],
     sp4_v_b_top[26], sp4_v_b_top[10], sp4_v_b_top[40],
     sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38], sp4_v_b_top[22],
     sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20], sp4_v_b_top[4],
     sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2], sp4_v_b_top[32],
     sp4_v_b_top[16], sp4_v_b_top[0]}), .sp4_r_v_b({sp4_r_v_b_top[47],
     sp4_r_v_b_top[31], sp4_r_v_b_top[15], sp4_r_v_b_top[45],
     sp4_r_v_b_top[29], sp4_r_v_b_top[13], sp4_r_v_b_top[43],
     sp4_r_v_b_top[27], sp4_r_v_b_top[11], sp4_r_v_b_top[41],
     sp4_r_v_b_top[25], sp4_r_v_b_top[9], sp4_r_v_b_top[39],
     sp4_r_v_b_top[23], sp4_r_v_b_top[7], sp4_r_v_b_top[37],
     sp4_r_v_b_top[21], sp4_r_v_b_top[5], sp4_r_v_b_top[35],
     sp4_r_v_b_top[19], sp4_r_v_b_top[3], sp4_r_v_b_top[33],
     sp4_r_v_b_top[17], sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46],
     sp4_h_r_top[30], sp4_h_r_top[14], sp4_h_r_top[44],
     sp4_h_r_top[28], sp4_h_r_top[12], sp4_h_r_top[42],
     sp4_h_r_top[26], sp4_h_r_top[10], sp4_h_r_top[40],
     sp4_h_r_top[24], sp4_h_r_top[8], sp4_h_r_top[38], sp4_h_r_top[22],
     sp4_h_r_top[6], sp4_h_r_top[36], sp4_h_r_top[20], sp4_h_r_top[4],
     sp4_h_r_top[34], sp4_h_r_top[18], sp4_h_r_top[2], sp4_h_r_top[32],
     sp4_h_r_top[16], sp4_h_r_top[0]}), .in3(bm_bweb[15:8]),
     .in2(in2_top[7:0]), .in1(bm_d[15:8]), .in0(net343[0:7]));

endmodule
// Library - leafcell, Cell - bram_4k_sr_bankout, View - schematic
// LAST TIME SAVED: Jul 25 22:59:22 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4k_sr_bankout ( bm_dm, bm_sdo, bm_sweb, clk, rcapmux_en,
     rst, bm_q, bm_sdi, wdummymux_en );
output  bm_sdo;

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[0]), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));
leafcell_ml_dff_schematic I29 ( .R(rst), .D(net0151), .CLK(clk),
     .QN(net0160), .Q(bm_sdo));
leafcell_ml_dff_schematic I22 ( .R(rst), .D(bm_dm[14]), .CLK(clk),
     .QN(net165), .Q(rdummy_reg));
ml_mux2_hvt_schematic I21 ( .in1(rdummy_reg), .in0(bm_dm[15]),
     .out(net0151), .sel(rdummymux_en));
nor2_hvt I24 ( .A(bm_swe), .B(rcapmux_en), .Y(net148));
inv_hvt I19 ( .A(bm_sweb), .Y(bm_swe));
inv_hvt I23 ( .A(net148), .Y(rdummymux_en));

endmodule
// Library - leafcell, Cell - bram_4k_bankout, View - schematic
// LAST TIME SAVED: Aug 15 18:09:39 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4k_bankout ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_ab;
input [7:0]  bm_sa;
input [7:0]  bm_aa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [15:0]  bm_dm;



tielo I15 ( .tielo(net092));
tielo I18 ( .tielo(net093));
bram_4k_sr_bankout I12 ( .bm_dm(bm_dm[15:0]), .rst(net093),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]), .bm_sdo(bm_sdo));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM(bm_dm[15:0]), .WEBM(bm_sweb), .WEB(web), .REBM(bm_sreb),
     .REB(reb), .D(bm_d[15:0]), .CLKW(net074), .CLKR(net072),
     .BWEBM({net092, net092, net092, net092, net092, net092, net092,
     net092, net092, net092, net092, net092, net092, net092, net092,
     net092}), .BWEB(bm_bweb[15:0]), .BIST(bm_init), .AMB(bm_sa[7:0]),
     .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]), .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net89), .out(net072));
bram_bufferx6 I8 ( .in(net85), .out(net074));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net85), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net89), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - leafcell, Cell - bram_4kbankout_pbuffer_bot, View -
//schematic
// LAST TIME SAVED: Aug 24 17:34:26 2007
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4kbankout_pbuffer_bot ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sdi_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sclkrw_o;

input [7:0]  bm_aa;
input [15:0]  bm_bweb;
input [7:0]  bm_sa_i;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sclkrw_i;
input [1:0]  bm_sdo_i;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [1:0]  bm_sweb_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o[0]), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i[0]), .bm_sclkrw_o(bm_sclkrw_o[0]),
     .bm_sdi_o(bm_sdi_o[0]), .bm_sdi_i(bm_sdi_i[0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k_bankout I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - misc, Cell - ml_osc_stage, View - schematic
// LAST TIME SAVED: Sep  8 19:15:04 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_osc_stage ( out, clkin, oscen_b, pbias, sel_trim );
output  out;

input  clkin, oscen_b, pbias;

input [3:0]  sel_trim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_mux3_hvt Iml_mux3_hvt_bot ( .in1(loadbot_1), .in0(loadbot_0),
     .out(in_bot), .sel(sel_trim[3:0]), .in2(loadbot_2));
nor2_hvt I228 ( .A(clkin), .B(oscen_b), .Y(net403));
inv_hvt I229 ( .A(net403), .Y(net419));
nch_hvt  MN41 ( .D(loadbot_0), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN39 ( .D(loadbot_2), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN29 ( .D(out), .B(gnd_), .G(in_bot), .S(gnd_));
nch_hvt  MN42 ( .D(loadbot_1), .B(gnd_), .G(net419), .S(gnd_));
pch_hvt  M82 ( .D(vdd_), .B(vdd_), .G(loadbot_1), .S(vdd_));
pch_hvt  M83 ( .D(vdd_), .B(vdd_), .G(loadbot_0), .S(vdd_));
pch_hvt  M85 ( .D(vdd_), .B(vdd_), .G(loadbot_2), .S(vdd_));
pch_hvt  M84 ( .D(vdd_), .B(vdd_), .G(loadbot_1), .S(vdd_));
pch_hvt  M81 ( .D(vdd_), .B(vdd_), .G(loadbot_2), .S(vdd_));
pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(loadbot_0), .S(vdd_));
pch_hvt  MP73 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net456));
pch_hvt  MP30 ( .D(net452), .B(vdd_), .G(oscen_b), .S(vdd_));
pch_hvt  MP72 ( .D(net456), .B(vdd_), .G(sel_trim[2]), .S(net452));
pch_hvt  MP33 ( .D(out), .B(vdd_), .G(in_bot), .S(vdd_));
pch_hvt  MP74 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net452));

endmodule
// Library - leafcell, Cell - bram_4kprouting_bbankout, View -
//schematic
// LAST TIME SAVED: Jan  8 10:35:21 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module bram_4kprouting_bbankout ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;
output [1:0]  bm_sclkrw_o;

inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_h_l_top;
inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_v_b_top;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_v_b_bot;
inout [23:0]  sp12_h_r_bot;
inout [47:0]  sp4_v_b_bot;
inout [41:0]  bl;
inout [47:0]  sp4_h_l_bot;

input [7:0]  top_op_top;
input [1:0]  bm_sclkrw_i;
input [1:0]  bm_sdi_i;
input [7:0]  glb_netwk;
input [7:0]  rgt_op_top;
input [7:0]  bnr_op_top;
input [7:0]  bot_op_bot;
input [7:0]  bm_sa_i;
input [7:0]  bnr_op_bot;
input [1:0]  bm_sdo_i;
input [15:0]  vdd_cntl_top;
input [7:0]  tnr_op_top;
input [7:0]  rgt_op_bot;
input [15:0]  wl_top;
input [15:0]  pgate_top;
input [15:0]  pgate_bot;
input [15:0]  reset_b_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  tnl_op_top;
input [1:0]  bm_sweb_i;
input [7:0]  bnl_op_top;
input [15:0]  reset_b_bot;
input [15:0]  wl_bot;
input [7:0]  lft_op_top;
input [7:0]  bnl_op_bot;
input [7:0]  tnl_op_bot;
input [7:0]  tnr_op_bot;
input [7:0]  lft_op_bot;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net252;

wire  [0:7]  net285;

wire  [0:7]  net341;

wire  [0:7]  net320;

wire  [7:0]  in2_top;

wire  [0:7]  net254;

wire  [0:7]  net286;

wire  [0:7]  net284;

wire  [0:7]  net253;

wire  [0:7]  net0239;

wire  [0:7]  net251;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net283;

wire  [15:0]  bm_d;

wire  [15:0]  bm_bweb;

wire  [0:7]  net0207;



bram_routing_tracks4rev12 I_bot ( .cbit_colcntl(net0207[0:7]),
     .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15], vdd_cntl_bot[12],
     vdd_cntl_bot[13], vdd_cntl_bot[10], vdd_cntl_bot[11],
     vdd_cntl_bot[8], vdd_cntl_bot[9], vdd_cntl_bot[6],
     vdd_cntl_bot[7], vdd_cntl_bot[4], vdd_cntl_bot[5],
     vdd_cntl_bot[2], vdd_cntl_bot[3], vdd_cntl_bot[0],
     vdd_cntl_bot[1]}), .s_r(net234), .wl({wl_bot[14], wl_bot[15],
     wl_bot[12], wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8],
     wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2],
     wl_bot[3], wl_bot[0], wl_bot[1]}), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net251[0:7]),
     .lc_trk_g2(net252[0:7]), .lc_trk_g1(net253[0:7]),
     .lc_trk_g0(net254[0:7]), .clk(net255),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev12 I_top ( .cbit_colcntl(net0239[0:7]),
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .s_r(net266), .wl({wl_top[14], wl_top[15],
     wl_top[12], wl_top[13], wl_top[10], wl_top[11], wl_top[8],
     wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2],
     wl_top[3], wl_top[0], wl_top[1]}), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net283[0:7]),
     .lc_trk_g2(net284[0:7]), .lc_trk_g1(net285[0:7]),
     .lc_trk_g0(net286[0:7]), .clk(net287),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbankout_pbuffer_bot I_bram_4kbankout_pbuffer_bot (
     .bm_q({slf_op_top[7:0], slf_op_bot[7:0]}),
     .bm_sdo_i(bm_sdo_i[1:0]), .bm_sdi_o(bm_sdi_o[1:0]),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sdi_i(bm_sdi_i[1:0]),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .bm_sweb_i(bm_sweb_i[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sweb_o(bm_sweb_o[1:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_init_i(bm_init_i),
     .bm_ren(net266), .bm_wen(net234), .bm_d(bm_d[15:0]),
     .bm_clkr(net287), .bm_clkw(net255), .bm_bweb(bm_bweb[15:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_ab(net341[0:7]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sreb_i(bm_sreb_i), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_aa(net320[0:7]), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_b ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}),
     .bl(bl[41:26]), .wl({wl_bot[14], wl_bot[15], wl_bot[12],
     wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8], wl_bot[9],
     wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2], wl_bot[3],
     wl_bot[0], wl_bot[1]}), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .op(slf_op_bot[7:0]), .lc_trk_g3(net251[0:7]),
     .lc_trk_g2(net252[0:7]), .lc_trk_g1(net253[0:7]),
     .lc_trk_g0(net254[0:7]), .sp12_h_r({sp12_h_r_bot[22],
     sp12_h_r_bot[6], sp12_h_r_bot[20], sp12_h_r_bot[4],
     sp12_h_r_bot[18], sp12_h_r_bot[2], sp12_h_r_bot[16],
     sp12_h_r_bot[0], sp12_h_r_bot[14], sp12_h_r_bot[12],
     sp12_h_r_bot[10], sp12_h_r_bot[8]}), .sp4_v_b({sp4_v_b_bot[46],
     sp4_v_b_bot[30], sp4_v_b_bot[14], sp4_v_b_bot[44],
     sp4_v_b_bot[28], sp4_v_b_bot[12], sp4_v_b_bot[42],
     sp4_v_b_bot[26], sp4_v_b_bot[10], sp4_v_b_bot[40],
     sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38], sp4_v_b_bot[22],
     sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20], sp4_v_b_bot[4],
     sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2], sp4_v_b_bot[32],
     sp4_v_b_bot[16], sp4_v_b_bot[0]}), .sp4_r_v_b({sp4_r_v_b_bot[47],
     sp4_r_v_b_bot[31], sp4_r_v_b_bot[15], sp4_r_v_b_bot[45],
     sp4_r_v_b_bot[29], sp4_r_v_b_bot[13], sp4_r_v_b_bot[43],
     sp4_r_v_b_bot[27], sp4_r_v_b_bot[11], sp4_r_v_b_bot[41],
     sp4_r_v_b_bot[25], sp4_r_v_b_bot[9], sp4_r_v_b_bot[39],
     sp4_r_v_b_bot[23], sp4_r_v_b_bot[7], sp4_r_v_b_bot[37],
     sp4_r_v_b_bot[21], sp4_r_v_b_bot[5], sp4_r_v_b_bot[35],
     sp4_r_v_b_bot[19], sp4_r_v_b_bot[3], sp4_r_v_b_bot[33],
     sp4_r_v_b_bot[17], sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46],
     sp4_h_r_bot[30], sp4_h_r_bot[14], sp4_h_r_bot[44],
     sp4_h_r_bot[28], sp4_h_r_bot[12], sp4_h_r_bot[42],
     sp4_h_r_bot[26], sp4_h_r_bot[10], sp4_h_r_bot[40],
     sp4_h_r_bot[24], sp4_h_r_bot[8], sp4_h_r_bot[38], sp4_h_r_bot[22],
     sp4_h_r_bot[6], sp4_h_r_bot[36], sp4_h_r_bot[20], sp4_h_r_bot[4],
     sp4_h_r_bot[34], sp4_h_r_bot[18], sp4_h_r_bot[2], sp4_h_r_bot[32],
     sp4_h_r_bot[16], sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]),
     .in2(in2_bot[7:0]), .in1(bm_d[7:0]), .in0(net320[0:7]),
     .sp12_v_b({sp12_v_b_bot[14], sp12_v_b_bot[12], sp12_v_b_bot[10],
     sp12_v_b_bot[8], sp12_v_b_bot[22], sp12_v_b_bot[6],
     sp12_v_b_bot[20], sp12_v_b_bot[4], sp12_v_b_bot[18],
     sp12_v_b_bot[2], sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_t ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}),
     .bl(bl[41:26]), .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12],
     sp12_v_b_top[10], sp12_v_b_top[8], sp12_v_b_top[22],
     sp12_v_b_top[6], sp12_v_b_top[20], sp12_v_b_top[4],
     sp12_v_b_top[18], sp12_v_b_top[2], sp12_v_b_top[16],
     sp12_v_b_top[0]}), .wl({wl_top[14], wl_top[15], wl_top[12],
     wl_top[13], wl_top[10], wl_top[11], wl_top[8], wl_top[9],
     wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2], wl_top[3],
     wl_top[0], wl_top[1]}), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .op(slf_op_top[7:0]), .lc_trk_g3(net283[0:7]),
     .lc_trk_g2(net284[0:7]), .lc_trk_g1(net285[0:7]),
     .lc_trk_g0(net286[0:7]), .sp12_h_r({sp12_h_r_top[22],
     sp12_h_r_top[6], sp12_h_r_top[20], sp12_h_r_top[4],
     sp12_h_r_top[18], sp12_h_r_top[2], sp12_h_r_top[16],
     sp12_h_r_top[0], sp12_h_r_top[14], sp12_h_r_top[12],
     sp12_h_r_top[10], sp12_h_r_top[8]}), .sp4_v_b({sp4_v_b_top[46],
     sp4_v_b_top[30], sp4_v_b_top[14], sp4_v_b_top[44],
     sp4_v_b_top[28], sp4_v_b_top[12], sp4_v_b_top[42],
     sp4_v_b_top[26], sp4_v_b_top[10], sp4_v_b_top[40],
     sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38], sp4_v_b_top[22],
     sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20], sp4_v_b_top[4],
     sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2], sp4_v_b_top[32],
     sp4_v_b_top[16], sp4_v_b_top[0]}), .sp4_r_v_b({sp4_r_v_b_top[47],
     sp4_r_v_b_top[31], sp4_r_v_b_top[15], sp4_r_v_b_top[45],
     sp4_r_v_b_top[29], sp4_r_v_b_top[13], sp4_r_v_b_top[43],
     sp4_r_v_b_top[27], sp4_r_v_b_top[11], sp4_r_v_b_top[41],
     sp4_r_v_b_top[25], sp4_r_v_b_top[9], sp4_r_v_b_top[39],
     sp4_r_v_b_top[23], sp4_r_v_b_top[7], sp4_r_v_b_top[37],
     sp4_r_v_b_top[21], sp4_r_v_b_top[5], sp4_r_v_b_top[35],
     sp4_r_v_b_top[19], sp4_r_v_b_top[3], sp4_r_v_b_top[33],
     sp4_r_v_b_top[17], sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46],
     sp4_h_r_top[30], sp4_h_r_top[14], sp4_h_r_top[44],
     sp4_h_r_top[28], sp4_h_r_top[12], sp4_h_r_top[42],
     sp4_h_r_top[26], sp4_h_r_top[10], sp4_h_r_top[40],
     sp4_h_r_top[24], sp4_h_r_top[8], sp4_h_r_top[38], sp4_h_r_top[22],
     sp4_h_r_top[6], sp4_h_r_top[36], sp4_h_r_top[20], sp4_h_r_top[4],
     sp4_h_r_top[34], sp4_h_r_top[18], sp4_h_r_top[2], sp4_h_r_top[32],
     sp4_h_r_top[16], sp4_h_r_top[0]}), .in3(bm_bweb[15:8]),
     .in2(in2_top[7:0]), .in1(bm_d[15:8]), .in0(net341[0:7]));

endmodule
// Library - leafcell, Cell - ice1f_array_BRAM_bot, View - schematic
// LAST TIME SAVED: Feb 12 17:38:41 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module ice1f_array_BRAM_bot ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, glb_netwk_bot, glb_netwk_top, slf_op_01,
     slf_op_02, slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07,
     slf_op_08, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02, sp4_h_l_03,
     sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07, sp4_h_l_08,
     sp4_h_r_01, sp4_h_r_02, sp4_h_r_03, sp4_h_r_04, sp4_h_r_05,
     sp4_h_r_06, sp4_h_r_07, sp4_h_r_08, sp4_r_v_b_01, sp4_r_v_b_02,
     sp4_r_v_b_03, sp4_r_v_b_04, sp4_r_v_b_05, sp4_r_v_b_06,
     sp4_r_v_b_07, sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03,
     sp4_v_b_04, sp4_v_b_05, sp4_v_b_06, sp4_v_b_07, sp4_v_b_08,
     sp4_v_t_08, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04,
     sp12_h_l_05, sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_r_01,
     sp12_h_r_02, sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06,
     sp12_h_r_07, sp12_h_r_08, sp12_v_b_01, sp12_v_t_08, vdd_cntl, wl,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i,
     bnl_op_01, bnr_op_01, bot_op_01, glb_netwk_col, lft_op_01,
     lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06, lft_op_07,
     lft_op_08, prog, rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04,
     rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, tnl_op_08, tnr_op_08,
     top_op_08 );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_05;
output [7:0]  slf_op_04;
output [1:0]  bm_sclkrw_o;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_07;
output [7:0]  slf_op_08;
output [7:0]  slf_op_01;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_03;
output [7:0]  slf_op_02;
output [7:0]  glb_netwk_bot;
output [7:0]  glb_netwk_top;
output [7:0]  slf_op_06;

inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_r_v_b_02;
inout [23:0]  sp12_h_l_01;
inout [23:0]  sp12_h_r_08;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_h_l_08;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_v_b_05;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_v_b_04;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_v_t_08;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_r_v_b_06;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_r_v_b_05;
inout [23:0]  sp12_v_t_08;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_h_l_02;
inout [23:0]  sp12_h_l_03;
inout [23:0]  sp12_h_l_07;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_h_r_03;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_r_v_b_04;
inout [47:0]  sp4_h_l_04;
inout [23:0]  sp12_h_l_04;
inout [47:0]  sp4_v_b_07;
inout [47:0]  sp4_v_b_08;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_h_l_03;
inout [47:0]  sp4_v_b_06;
inout [47:0]  sp4_h_l_01;
inout [47:0]  sp4_v_b_03;
inout [23:0]  sp12_h_r_04;
inout [127:0]  wl;
inout [127:0]  vdd_cntl;
inout [127:0]  reset_b;
inout [127:0]  pgate;
inout [47:0]  sp4_h_r_08;
inout [47:0]  sp4_h_r_04;
inout [23:0]  sp12_h_l_06;
inout [41:0]  bl;
inout [47:0]  sp4_h_l_07;
inout [47:0]  sp4_r_v_b_01;
inout [23:0]  sp12_v_b_01;
inout [47:0]  sp4_h_l_06;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_h_l_05;
inout [23:0]  sp12_h_l_05;
inout [23:0]  sp12_h_r_06;

input [7:0]  rgt_op_01;
input [7:0]  rgt_op_04;
input [7:0]  lft_op_02;
input [7:0]  tnl_op_08;
input [1:0]  bm_sclkrw_i;
input [7:0]  rgt_op_07;
input [1:0]  bm_sweb_i;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_03;
input [7:0]  rgt_op_08;
input [7:0]  lft_op_01;
input [7:0]  rgt_op_06;
input [7:0]  bnl_op_01;
input [1:0]  bm_sdi_i;
input [7:0]  top_op_08;
input [7:0]  lft_op_06;
input [7:0]  lft_op_08;
input [1:0]  bm_sdo_i;
input [7:0]  bot_op_01;
input [7:0]  bnr_op_01;
input [7:0]  lft_op_04;
input [7:0]  glb_netwk_col;
input [7:0]  lft_op_07;
input [7:0]  lft_op_05;
input [7:0]  tnr_op_08;
input [7:0]  bm_sa_i;
input [7:0]  rgt_op_02;
input [7:0]  lft_op_03;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  colbuf_cntl_bot;

wire  [7:0]  colbuf_cntl_top;

wire  [0:7]  net0808;

wire  [0:1]  net0863;

wire  [0:1]  net0862;

wire  [0:23]  net1169;

wire  [0:1]  net0866;

wire  [0:23]  net1107;

wire  [0:7]  net1133;

wire  [0:1]  net0930;

wire  [0:1]  net0868;

wire  [0:7]  net823;

wire  [0:1]  net01362;

wire  [0:1]  net01359;

wire  [0:1]  net01358;

wire  [0:1]  net0928;

wire  [0:7]  net1195;

wire  [0:1]  net0924;

wire  [0:23]  net797;

wire  [0:1]  net01364;

wire  [0:1]  net0925;



clk_colbuf1kx8 I_clk_colbuf12kx8_b (
     .colbuf_cntl(colbuf_cntl_bot[7:0]), .col_clk(glb_netwk_bot[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_colbuf1kx8 I_clk_colbuf12kx8_t (
     .colbuf_cntl(colbuf_cntl_top[7:0]), .col_clk(glb_netwk_top[7:0]),
     .clk_in(glb_netwk_col[7:0]));
bram_4kprouting_bbank I_bram_0708 ( .cbit_colcntl(net0808[0:7]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sclkrw_i(net0925[0:1]), .bm_sweb_i(net0928[0:1]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_sdi_i(net0924[0:1]),
     .bm_sdo_i(bm_sdo_i[1:0]), .bm_sdo_o(net0930[0:1]),
     .slf_op_top(slf_op_08[7:0]), .slf_op_bot(slf_op_07[7:0]),
     .wl_bot(wl[111:96]), .top_op_top(top_op_08[7:0]),
     .sp12_h_l_bot(sp12_h_l_07[23:0]), .sp4_h_l_bot(sp4_h_l_07[47:0]),
     .tnl_op_top(tnl_op_08[7:0]), .tnl_op_bot(lft_op_08[7:0]),
     .reset_b_top(reset_b[127:112]), .reset_b_bot(reset_b[111:96]),
     .vdd_cntl_top(vdd_cntl[127:112]), .prog(prog),
     .pgate_top(pgate[127:112]), .pgate_bot(pgate[111:96]),
     .lft_op_bot(lft_op_07[7:0]), .glb_netwk(glb_netwk_top[7:0]),
     .bm_wdummymux_en_i(net1136), .bot_op_bot(slf_op_06[7:0]),
     .rgt_op_bot(rgt_op_07[7:0]), .bnl_op_top(lft_op_07[7:0]),
     .bnl_op_bot(lft_op_06[7:0]), .sp4_h_r_top(sp4_h_r_08[47:0]),
     .sp12_v_t_top(sp12_v_t_08[23:0]), .sp12_v_b_bot(net1107[0:23]),
     .bm_init_i(net1132), .sp4_h_r_bot(sp4_h_r_07[47:0]),
     .sp12_h_r_bot(sp12_h_r_07[23:0]), .sp4_v_t_top(sp4_v_t_08[47:0]),
     .sp4_v_b_bot(sp4_v_b_07[47:0]), .sp12_h_r_top(sp12_h_r_08[23:0]),
     .tnr_op_bot(rgt_op_08[7:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(net1131), .sp4_h_l_top(sp4_h_l_08[47:0]),
     .lft_op_top(lft_op_08[7:0]), .wl_top(wl[127:112]),
     .sp12_h_l_top(sp12_h_l_08[23:0]), .sp4_v_b_top(sp4_v_b_08[47:0]),
     .tnr_op_top(tnr_op_08[7:0]), .rgt_op_top(rgt_op_08[7:0]),
     .bm_sa_i(net1133[0:7]), .bm_sclk_i(net1134), .bm_sreb_i(net1135),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .vdd_cntl_bot(vdd_cntl[111:96]), .bnr_op_bot(rgt_op_06[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_07[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_08[47:0]), .bnr_op_top(rgt_op_07[7:0]));
bram_4kprouting_bbank I_bram_0506 (
     .cbit_colcntl(colbuf_cntl_top[7:0]), .bm_sdi_o(net0924[0:1]),
     .bm_sclkrw_o(net0925[0:1]), .bm_sclkrw_i(net0863[0:1]),
     .bm_sweb_i(net0866[0:1]), .bm_sweb_o(net0928[0:1]),
     .bm_sdi_i(net0862[0:1]), .bm_sdo_i(net0930[0:1]),
     .bm_sdo_o(net0868[0:1]), .slf_op_top(slf_op_06[7:0]),
     .slf_op_bot(slf_op_05[7:0]), .wl_top(wl[95:80]),
     .wl_bot(wl[79:64]), .top_op_top(slf_op_07[7:0]),
     .tnl_op_top(lft_op_07[7:0]), .tnl_op_bot(lft_op_06[7:0]),
     .reset_b_top(reset_b[95:80]), .reset_b_bot(reset_b[79:64]),
     .prog(prog), .pgate_top(pgate[95:80]), .pgate_bot(pgate[79:64]),
     .lft_op_top(lft_op_06[7:0]), .lft_op_bot(lft_op_05[7:0]),
     .glb_netwk(glb_netwk_top[7:0]), .bm_wdummymux_en_i(net1198),
     .bot_op_bot(slf_op_04[7:0]), .sp4_h_r_top(sp4_h_r_06[47:0]),
     .bnl_op_top(lft_op_05[7:0]), .bnl_op_bot(lft_op_04[7:0]),
     .bnr_op_bot(rgt_op_04[7:0]), .sp4_h_r_bot(sp4_h_r_05[47:0]),
     .sp12_v_t_top(net1107[0:23]), .sp12_v_b_bot(net1169[0:23]),
     .bm_init_i(net1194), .sp12_h_l_top(sp12_h_l_06[23:0]),
     .sp12_h_r_bot(sp12_h_r_05[23:0]),
     .sp12_h_l_bot(sp12_h_l_05[23:0]),
     .sp12_h_r_top(sp12_h_r_06[23:0]), .sp4_v_t_top(sp4_v_b_07[47:0]),
     .sp4_v_b_top(sp4_v_b_06[47:0]), .sp4_v_b_bot(sp4_v_b_05[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_05[47:0]),
     .sp4_h_l_top(sp4_h_l_06[47:0]), .tnr_op_top(rgt_op_07[7:0]),
     .sp4_h_l_bot(sp4_h_l_05[47:0]), .tnr_op_bot(rgt_op_06[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net1193),
     .sp4_r_v_b_top(sp4_r_v_b_06[47:0]), .rgt_op_bot(rgt_op_05[7:0]),
     .rgt_op_top(rgt_op_06[7:0]), .bnr_op_top(rgt_op_05[7:0]),
     .bm_sa_i(net1195[0:7]), .bm_sclk_i(net1196), .bm_sreb_i(net1197),
     .bm_rcapmux_en_o(net1131), .bm_init_o(net1132),
     .bm_sa_o(net1133[0:7]), .bm_sclk_o(net1134), .bm_sreb_o(net1135),
     .bm_wdummymux_en_o(net1136), .vdd_cntl_top(vdd_cntl[95:80]),
     .vdd_cntl_bot(vdd_cntl[79:64]));
bram_4kprouting_bbank I_bram_0304 (
     .cbit_colcntl(colbuf_cntl_bot[7:0]), .bm_sdi_o(net0862[0:1]),
     .bm_sclkrw_o(net0863[0:1]), .bm_sclkrw_i(net01359[0:1]),
     .bm_sweb_i(net01362[0:1]), .bm_sweb_o(net0866[0:1]),
     .bm_sdi_i(net01358[0:1]), .bm_sdo_i(net0868[0:1]),
     .bm_sdo_o(net01364[0:1]), .slf_op_top(slf_op_04[7:0]),
     .slf_op_bot(slf_op_03[7:0]), .wl_top(wl[63:48]),
     .wl_bot(wl[47:32]), .top_op_top(slf_op_05[7:0]),
     .tnl_op_top(lft_op_05[7:0]), .tnl_op_bot(lft_op_04[7:0]),
     .reset_b_top(reset_b[63:48]), .reset_b_bot(reset_b[47:32]),
     .prog(prog), .pgate_top(pgate[63:48]), .pgate_bot(pgate[47:32]),
     .lft_op_top(lft_op_04[7:0]), .lft_op_bot(lft_op_03[7:0]),
     .glb_netwk(glb_netwk_bot[7:0]), .bm_wdummymux_en_i(net826),
     .bot_op_bot(slf_op_02[7:0]), .sp4_h_r_top(sp4_h_r_04[47:0]),
     .bnl_op_top(lft_op_03[7:0]), .bnl_op_bot(lft_op_02[7:0]),
     .bnr_op_bot(rgt_op_02[7:0]), .sp4_h_r_bot(sp4_h_r_03[47:0]),
     .sp12_v_t_top(net1169[0:23]), .sp12_v_b_bot(net797[0:23]),
     .bm_init_i(net822), .sp12_h_l_top(sp12_h_l_04[23:0]),
     .sp12_h_r_bot(sp12_h_r_03[23:0]),
     .sp12_h_l_bot(sp12_h_l_03[23:0]),
     .sp12_h_r_top(sp12_h_r_04[23:0]), .sp4_v_t_top(sp4_v_b_05[47:0]),
     .sp4_v_b_top(sp4_v_b_04[47:0]), .sp4_v_b_bot(sp4_v_b_03[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_03[47:0]),
     .sp4_h_l_top(sp4_h_l_04[47:0]), .tnr_op_top(rgt_op_05[7:0]),
     .sp4_h_l_bot(sp4_h_l_03[47:0]), .tnr_op_bot(rgt_op_04[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net821),
     .sp4_r_v_b_top(sp4_r_v_b_04[47:0]), .rgt_op_bot(rgt_op_03[7:0]),
     .rgt_op_top(rgt_op_04[7:0]), .bnr_op_top(rgt_op_03[7:0]),
     .bm_sa_i(net823[0:7]), .bm_sclk_i(net824), .bm_sreb_i(net825),
     .bm_rcapmux_en_o(net1193), .bm_init_o(net1194),
     .bm_sa_o(net1195[0:7]), .bm_sclk_o(net1196), .bm_sreb_o(net1197),
     .bm_wdummymux_en_o(net1198), .vdd_cntl_top(vdd_cntl[63:48]),
     .vdd_cntl_bot(vdd_cntl[47:32]));
bram_4kprouting_bbankout I_bram_out_0102 ( .bm_sdi_o(net01358[0:1]),
     .bm_sclkrw_o(net01359[0:1]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sweb_o(net01362[0:1]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sdo_i(net01364[0:1]),
     .bm_sdo_o(bm_sdo_o[1:0]), .slf_op_top(slf_op_02[7:0]),
     .slf_op_bot(slf_op_01[7:0]), .wl_top(wl[31:16]),
     .wl_bot(wl[15:0]), .top_op_top(slf_op_03[7:0]),
     .tnl_op_top(lft_op_03[7:0]), .tnl_op_bot(lft_op_02[7:0]),
     .reset_b_top(reset_b[31:16]), .reset_b_bot(reset_b[15:0]),
     .prog(prog), .pgate_top(pgate[31:16]), .pgate_bot(pgate[15:0]),
     .lft_op_top(lft_op_02[7:0]), .lft_op_bot(lft_op_01[7:0]),
     .glb_netwk(glb_netwk_bot[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bot_op_bot(bot_op_01[7:0]), .sp4_h_r_top(sp4_h_r_02[47:0]),
     .bnl_op_top(lft_op_01[7:0]), .bnl_op_bot(bnl_op_01[7:0]),
     .bnr_op_bot(bnr_op_01[7:0]), .sp4_h_r_bot(sp4_h_r_01[47:0]),
     .sp12_v_t_top(net797[0:23]), .sp12_v_b_bot(sp12_v_b_01[23:0]),
     .bm_init_i(bm_init_i), .sp12_h_l_top(sp12_h_l_02[23:0]),
     .sp12_h_r_bot(sp12_h_r_01[23:0]),
     .sp12_h_l_bot(sp12_h_l_01[23:0]),
     .sp12_h_r_top(sp12_h_r_02[23:0]), .sp4_v_t_top(sp4_v_b_03[47:0]),
     .sp4_v_b_top(sp4_v_b_02[47:0]), .sp4_v_b_bot(sp4_v_b_01[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_01[47:0]),
     .sp4_h_l_top(sp4_h_l_02[47:0]), .tnr_op_top(rgt_op_03[7:0]),
     .sp4_h_l_bot(sp4_h_l_01[47:0]), .tnr_op_bot(rgt_op_02[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .sp4_r_v_b_top(sp4_r_v_b_02[47:0]), .rgt_op_bot(rgt_op_01[7:0]),
     .rgt_op_top(rgt_op_02[7:0]), .bnr_op_top(rgt_op_01[7:0]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sreb_i(bm_sreb_i), .bm_rcapmux_en_o(net821),
     .bm_init_o(net822), .bm_sa_o(net823[0:7]), .bm_sclk_o(net824),
     .bm_sreb_o(net825), .bm_wdummymux_en_o(net826),
     .vdd_cntl_top(vdd_cntl[31:16]), .vdd_cntl_bot(vdd_cntl[15:0]));

endmodule
// Library - leafcell, Cell - fabric_outbuf12p, View - schematic
// LAST TIME SAVED: Dec 17 09:43:15 2008
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module fabric_outbuf12p ( cout, fabric_out );
output  cout;

input  fabric_out;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I24 ( .A(fabric_out), .Y(net19));
inv_hvt I23 ( .A(net19), .Y(cout));

endmodule
// Library - leafcell, Cell - clk_quadbuf12k, View - schematic
// LAST TIME SAVED: Mar 19 09:33:13 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module clk_quadbuf12k ( clko, clki );
output  clko;

input  clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I23 ( .A(clki), .Y(clkb));
inv_hvt I25 ( .A(clkb), .Y(clko));

endmodule
// Library - leafcell, Cell - clk_quad_buf12px8, View - schematic
// LAST TIME SAVED: Jan 21 11:21:33 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module clk_quad_buf12px8 ( clko, clki );


output [7:0]  clko;

input [7:0]  clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clk_quadbuf12k Iclk_quadbuf12k_7_ ( .clki(clki[7]), .clko(clko[7]));
clk_quadbuf12k Iclk_quadbuf12k_6_ ( .clki(clki[6]), .clko(clko[6]));
clk_quadbuf12k Iclk_quadbuf12k_5_ ( .clki(clki[5]), .clko(clko[5]));
clk_quadbuf12k Iclk_quadbuf12k_4_ ( .clki(clki[4]), .clko(clko[4]));
clk_quadbuf12k Iclk_quadbuf12k_3_ ( .clki(clki[3]), .clko(clko[3]));
clk_quadbuf12k Iclk_quadbuf12k_2_ ( .clki(clki[2]), .clko(clko[2]));
clk_quadbuf12k Iclk_quadbuf12k_1_ ( .clki(clki[1]), .clko(clko[1]));
clk_quadbuf12k Iclk_quadbuf12k_0_ ( .clki(clki[0]), .clko(clko[0]));

endmodule
// Library - leafcell, Cell - ice1f_quad_bl, View - schematic
// LAST TIME SAVED: Jul 22 09:11:58 2009
// NETLIST TIME: Aug 24 09:59:01 2009
`timescale 1ns / 1ns 

module ice1f_quad_bl ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_01_08, carry_out_02_08,
     carry_out_04_08, carry_out_05_08, carry_out_06_08, ceb_o, cf_b_l,
     cf_l, fabric_out_00_07, fabric_out_00_08, fabric_out_05_00,
     fabric_out_06_00, hiz_b_o, mode_o, padeb_b_l, padeb_l_b,
     padin_00_08b, padin_06_00b, pado_b_l, pado_l_b, r_o, sdo, shift_o,
     slf_op_00_08, slf_op_01_08, slf_op_02_08, slf_op_03_08,
     slf_op_04_08, slf_op_05_08, slf_op_06_00, slf_op_06_01,
     slf_op_06_02, slf_op_06_03, slf_op_06_04, slf_op_06_05,
     slf_op_06_06, slf_op_06_07, slf_op_06_08, spi_ss_in_l, tclk_o,
     update_o, bl, pgate_l, reset_b_l, sp4_h_r_06_00, sp4_h_r_06_01,
     sp4_h_r_06_02, sp4_h_r_06_03, sp4_h_r_06_04, sp4_h_r_06_05,
     sp4_h_r_06_06, sp4_h_r_06_07, sp4_h_r_06_08, sp4_r_v_b_06_01,
     sp4_r_v_b_06_02, sp4_r_v_b_06_03, sp4_r_v_b_06_04,
     sp4_r_v_b_06_05, sp4_r_v_b_06_06, sp4_r_v_b_06_07,
     sp4_r_v_b_06_08, sp4_v_t_00_08, sp4_v_t_01_08, sp4_v_t_02_08,
     sp4_v_t_03_08, sp4_v_t_04_08, sp4_v_t_05_08, sp4_v_t_06_08,
     sp12_h_r_06_01, sp12_h_r_06_02, sp12_h_r_06_03, sp12_h_r_06_04,
     sp12_h_r_06_05, sp12_h_r_06_06, sp12_h_r_06_07, sp12_h_r_06_08,
     sp12_v_t_01_08, sp12_v_t_02_08, sp12_v_t_03_08, sp12_v_t_04_08,
     sp12_v_t_05_08, sp12_v_t_06_08, vdd_cntl_l, wl_l, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnr_op_06_01,
     bs_en_i, ceb_i, end_of_startup_lft_b, glb_in, hiz_b_i, hold_b_l,
     hold_l_b, mode_i, padin_b_l, padin_l_b, prog, purst, r_i,
     rgt_op_06_01, rgt_op_06_02, rgt_op_06_03, rgt_op_06_04,
     rgt_op_06_05, rgt_op_06_06, rgt_op_06_07, rgt_op_06_08, sdi,
     shift_i, spioeb_l, spiout_l, tclk_i, tiegnd, tievdd, tnl_op_01_08,
     tnl_op_02_08, tnl_op_03_08, tnl_op_04_08, tnl_op_05_08,
     tnl_op_06_08, tnr_op_00_08, tnr_op_01_08, tnr_op_02_08,
     tnr_op_03_08, tnr_op_04_08, tnr_op_05_08, tnr_op_06_00,
     tnr_op_06_08, top_op_01_08, top_op_02_08, top_op_03_08,
     top_op_04_08, top_op_05_08, top_op_06_08, update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_01_08, carry_out_02_08,
     carry_out_04_08, carry_out_05_08, carry_out_06_08, ceb_o,
     fabric_out_00_07, fabric_out_00_08, fabric_out_05_00,
     fabric_out_06_00, hiz_b_o, mode_o, padin_00_08b, padin_06_00b,
     r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, ceb_i, hiz_b_i, hold_b_l, hold_l_b,
     mode_i, prog, purst, r_i, sdi, shift_i, tclk_i, tiegnd, tievdd,
     update_i;

output [7:0]  slf_op_06_07;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_06_08;
output [7:0]  slf_op_06_05;
output [13:0]  pado_l_b;
output [7:0]  slf_op_05_08;
output [1:0]  bm_sclkrw_o;
output [3:0]  slf_op_00_08;
output [7:0]  slf_op_06_01;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_03_08;
output [7:0]  slf_op_06_03;
output [7:0]  slf_op_01_08;
output [7:0]  slf_op_06_04;
output [7:0]  slf_op_06_06;
output [13:0]  padeb_l_b;
output [7:0]  slf_op_04_08;
output [1:0]  bm_sdo_o;
output [15:0]  spi_ss_in_l;
output [11:0]  padeb_b_l;
output [143:0]  cf_b_l;
output [11:0]  pado_b_l;
output [191:0]  cf_l;
output [7:0]  slf_op_02_08;
output [7:0]  slf_op_06_02;
output [3:0]  slf_op_06_00;
output [7:0]  bm_sa_o;

inout [47:0]  sp4_r_v_b_06_07;
inout [23:0]  sp12_h_r_06_02;
inout [47:0]  sp4_h_r_06_01;
inout [23:0]  sp12_h_r_06_03;
inout [47:0]  sp4_h_r_06_05;
inout [47:0]  sp4_r_v_b_06_05;
inout [47:0]  sp4_v_t_03_08;
inout [47:0]  sp4_h_r_06_04;
inout [23:0]  sp12_h_r_06_05;
inout [47:0]  sp4_r_v_b_06_03;
inout [47:0]  sp4_r_v_b_06_08;
inout [23:0]  sp12_h_r_06_01;
inout [47:0]  sp4_h_r_06_07;
inout [47:0]  sp4_r_v_b_06_04;
inout [15:0]  sp4_v_t_00_08;
inout [23:0]  sp12_v_t_02_08;
inout [47:0]  sp4_h_r_06_06;
inout [47:0]  sp4_h_r_06_08;
inout [47:0]  sp4_v_t_01_08;
inout [23:0]  sp12_h_r_06_08;
inout [23:0]  sp12_h_r_06_04;
inout [47:0]  sp4_h_r_06_03;
inout [23:0]  sp12_v_t_04_08;
inout [23:0]  sp12_v_t_06_08;
inout [47:0]  sp4_r_v_b_06_01;
inout [47:0]  sp4_r_v_b_06_02;
inout [23:0]  sp12_v_t_03_08;
inout [23:0]  sp12_v_t_05_08;
inout [23:0]  sp12_h_r_06_06;
inout [47:0]  sp4_v_t_06_08;
inout [15:0]  sp4_h_r_06_00;
inout [47:0]  sp4_v_t_04_08;
inout [47:0]  sp4_v_t_05_08;
inout [23:0]  sp12_h_r_06_07;
inout [23:0]  sp12_v_t_01_08;
inout [143:0]  pgate_l;
inout [47:0]  sp4_r_v_b_06_06;
inout [47:0]  sp4_v_t_02_08;
inout [143:0]  reset_b_l;
inout [143:0]  vdd_cntl_l;
inout [329:0]  bl;
inout [143:0]  wl_l;
inout [47:0]  sp4_h_r_06_02;

input [7:0]  tnr_op_02_08;
input [7:0]  top_op_01_08;
input [7:0]  tnr_op_03_08;
input [7:0]  top_op_05_08;
input [7:0]  tnl_op_01_08;
input [13:0]  padin_l_b;
input [1:0]  bm_sclkrw_i;
input [7:0]  tnl_op_02_08;
input [1:0]  bm_sdi_i;
input [7:0]  rgt_op_06_08;
input [11:0]  padin_b_l;
input [7:0]  rgt_op_06_04;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_06_08;
input [7:0]  top_op_04_08;
input [3:0]  bnr_op_06_01;
input [7:0]  tnl_op_03_08;
input [7:0]  tnl_op_04_08;
input [7:0]  tnr_op_06_08;
input [7:0]  rgt_op_06_06;
input [7:0]  top_op_02_08;
input [7:0]  top_op_06_08;
input [7:0]  rgt_op_06_02;
input [15:0]  spioeb_l;
input [7:0]  tnr_op_05_08;
input [1:0]  bm_sdo_i;
input [7:0]  rgt_op_06_05;
input [7:0]  tnr_op_06_00;
input [7:0]  rgt_op_06_01;
input [7:0]  tnr_op_01_08;
input [7:0]  tnr_op_04_08;
input [8:1]  end_of_startup_lft_b;
input [7:0]  tnr_op_00_08;
input [1:0]  bm_sweb_i;
input [7:0]  tnl_op_05_08;
input [15:0]  spiout_l;
input [7:0]  rgt_op_06_03;
input [7:0]  top_op_03_08;
input [7:0]  rgt_op_06_07;
input [7:0]  glb_in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net1321;

wire  [0:23]  net1266;

wire  [0:7]  net837;

wire  [0:47]  net829;

wire  [0:23]  net1033;

wire  [0:23]  net1378;

wire  [0:47]  net831;

wire  [0:47]  net1381;

wire  [0:47]  net1134;

wire  [0:47]  net996;

wire  [0:7]  net1364;

wire  [0:47]  net1088;

wire  [0:47]  net1107;

wire  [0:47]  net1016;

wire  [0:7]  net731;

wire  [0:47]  net1137;

wire  [0:23]  net1171;

wire  [0:47]  net810;

wire  [0:23]  net1267;

wire  [0:47]  net1361;

wire  [0:47]  net1041;

wire  [0:47]  net1084;

wire  [0:47]  net1330;

wire  [0:47]  net686;

wire  [0:47]  net807;

wire  [0:47]  net1283;

wire  [0:47]  net1202;

wire  [0:23]  net1306;

wire  [0:47]  net990;

wire  [0:47]  net855;

wire  [0:23]  net1035;

wire  [0:47]  net1243;

wire  [0:47]  net1017;

wire  [0:47]  net1177;

wire  [0:23]  net798;

wire  [0:23]  net1366;

wire  [0:23]  net1129;

wire  [0:47]  net853;

wire  [0:7]  net1471;

wire  [0:7]  net1067;

wire  [0:23]  net849;

wire  [0:23]  net1172;

wire  [0:47]  net1175;

wire  [0:23]  net1221;

wire  [0:47]  net852;

wire  [0:7]  net1472;

wire  [0:47]  net690;

wire  [0:23]  net1076;

wire  [0:23]  net848;

wire  [0:47]  net1286;

wire  [0:47]  net1087;

wire  [0:23]  net705;

wire  [0:23]  net847;

wire  [0:23]  net1358;

wire  [0:47]  net698;

wire  [0:7]  net1437;

wire  [0:23]  net1305;

wire  [0:7]  net974;

wire  [0:47]  net1082;

wire  [0:7]  net966;

wire  [0:47]  net1014;

wire  [0:47]  net1373;

wire  [0:7]  net1384;

wire  [0:7]  net1057;

wire  [0:47]  net1181;

wire  [0:47]  net1333;

wire  [0:7]  net1435;

wire  [0:47]  net1279;

wire  [0:7]  net964;

wire  [0:23]  net799;

wire  [0:23]  net1362;

wire  [0:23]  net1370;

wire  [0:23]  net1382;

wire  [0:47]  net805;

wire  [0:47]  net1179;

wire  [0:47]  net1284;

wire  [0:7]  net1328;

wire  [0:47]  net1385;

wire  [0:47]  net1136;

wire  [0:7]  net1024;

wire  [0:47]  net994;

wire  [0:23]  net850;

wire  [0:23]  net800;

wire  [0:7]  net696;

wire  [0:7]  net1116;

wire  [0:47]  net1132;

wire  [0:7]  net1025;

wire  [0:23]  net1079;

wire  [0:7]  net1372;

wire  [0:7]  net1023;

wire  [0:23]  net1220;

wire  [0:47]  net854;

wire  [0:7]  net1315;

wire  [0:7]  net1452;

wire  [0:7]  net839;

wire  [0:23]  net697;

wire  [0:47]  net828;

wire  [0:7]  net1117;

wire  [0:47]  net1015;

wire  [0:47]  net1131;

wire  [0:7]  net788;

wire  [0:7]  net729;

wire  [0:7]  net838;

wire  [0:47]  net995;

wire  [0:23]  net1219;

wire  [0:23]  net983;

wire  [0:47]  net1039;

wire  [0:47]  net706;

wire  [0:47]  net1038;

wire  [3:0]  slf_op_00_03;

wire  [3:0]  slf_op_02_00;

wire  [0:47]  net702;

wire  [0:47]  net1099;

wire  [0:23]  net1036;

wire  [0:47]  net1133;

wire  [0:47]  net1180;

wire  [0:23]  net986;

wire  [0:47]  net1138;

wire  [0:47]  net1466;

wire  [0:23]  net1127;

wire  [0:23]  net701;

wire  [0:47]  net830;

wire  [0:7]  net726;

wire  [0:47]  net1303;

wire  [0:23]  net985;

wire  [0:23]  net1169;

wire  [0:23]  net1265;

wire  [13:13]  padinlat_l_b;

wire  [0:47]  net1110;

wire  [0:47]  net1086;

wire  [0:47]  net694;

wire  [0:47]  net803;

wire  [0:47]  net804;

wire  [0:23]  net1374;

wire  [3:0]  slf_op_05_00;

wire  [0:7]  net780;

wire  [3:0]  slf_op_00_01;

wire  [0:47]  net1331;

wire  [0:47]  net1340;

wire  [0:47]  net1338;

wire  [11:11]  padinlat_b_l;

wire  [0:7]  net1380;

wire  [0:47]  net1301;

wire  [0:23]  net1263;

wire  [3:0]  slf_op_00_06;

wire  [0:23]  net984;

wire  [0:23]  net1128;

wire  [0:47]  net1108;

wire  [0:23]  net709;

wire  [0:47]  net1365;

wire  [0:7]  net727;

wire  [0:47]  net1135;

wire  [0:47]  net1227;

wire  [3:0]  slf_op_01_00;

wire  [3:0]  slf_op_03_00;

wire  [0:47]  net808;

wire  [0:23]  net693;

wire  [0:47]  net1332;

wire  [3:0]  slf_op_00_07;

wire  [0:47]  net809;

wire  [0:47]  net1040;

wire  [0:47]  net1203;

wire  [3:0]  slf_op_00_02;

wire  [0:47]  net1101;

wire  [0:47]  net1109;

wire  [0:47]  net1201;

wire  [0:47]  net1100;

wire  [0:7]  net704;

wire  [0:23]  net1270;

wire  [0:47]  net1224;

wire  [0:7]  net1368;

wire  [0:23]  net797;

wire  [0:7]  net1318;

wire  [0:7]  net1319;

wire  [0:15]  net1397;

wire  [0:23]  net1308;

wire  [0:47]  net1226;

wire  [0:7]  net778;

wire  [0:47]  net989;

wire  [0:7]  net1059;

wire  [0:47]  net1176;

wire  [0:7]  net728;

wire  [0:7]  net1118;

wire  [0:7]  net1376;

wire  [0:47]  net993;

wire  [0:23]  net1034;

wire  [0:47]  net1089;

wire  [0:47]  net1083;

wire  [3:0]  slf_op_00_05;

wire  [0:7]  net730;

wire  [0:23]  net1386;

wire  [0:23]  net1078;

wire  [0:47]  net1225;

wire  [0:23]  net1077;

wire  [0:47]  net1369;

wire  [0:23]  net689;

wire  [0:7]  net1428;

wire  [0:7]  net692;

wire  [0:7]  net768;

wire  [0:47]  net1182;

wire  [0:23]  net1170;

wire  [0:7]  net1327;

wire  [0:47]  net1281;

wire  [0:23]  net1222;

wire  [3:0]  slf_op_04_00;

wire  [0:47]  net1377;

wire  [0:47]  net991;

wire  [0:47]  net1200;

wire  [3:0]  slf_op_00_04;

wire  [0:23]  net1126;

wire  [0:7]  net1453;

wire  [7:0]  clk_tree_drv;

wire  [0:47]  net1302;



ice1f_array_LFT_IO_bot14io I_preio_lft_b00 ( .padin(padin_l_b[13:0]),
     .pado(pado_l_b[13:0]), .padeb(padeb_l_b[13:0]),
     .sp4_v_t_00_08(sp4_v_t_00_08[15:0]),
     .tnl_op_00_08(tnr_op_00_08[7:0]),
     .cdone_in(end_of_startup_lft_b[8:1]), .wl(wl_l[143:16]),
     .vdd_cntl(vdd_cntl_l[143:16]), .reset_b(reset_b_l[143:16]),
     .pgate(pgate_l[143:16]), .spi_ss_in_b(spi_ss_in_l[15:0]),
     .spioeb(spioeb_l[15:0]), .spiout(spiout_l[15:0]),
     .cf_l(cf_l[191:0]), .bnl_op_00_01({slf_op_01_00[3],
     slf_op_01_00[2], slf_op_01_00[1], slf_op_01_00[0],
     slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0]}), .SP4_h_l_00_01(net1466[0:47]),
     .SP12_h_l_00_01(net1358[0:23]), .slf_op_00_01(slf_op_00_01[3:0]),
     .rgt_op_00_01(net1472[0:7]), .SP4_h_l_00_02(net1361[0:47]),
     .SP12_h_l_00_02(net1362[0:23]), .slf_op_00_02(slf_op_00_02[3:0]),
     .rgt_op_00_02(net1364[0:7]), .SP4_h_l_00_03(net1365[0:47]),
     .SP12_h_l_00_03(net1366[0:23]), .slf_op_00_03(slf_op_00_03[3:0]),
     .rgt_op_00_03(net1368[0:7]), .SP4_h_l_00_04(net1369[0:47]),
     .SP12_h_l_00_04(net1370[0:23]), .slf_op_00_04(slf_op_00_04[3:0]),
     .rgt_op_00_04(net1372[0:7]), .SP4_h_l_00_05(net1373[0:47]),
     .SP12_h_l_00_05(net1374[0:23]), .slf_op_00_05(slf_op_00_05[3:0]),
     .rgt_op_00_05(net1376[0:7]), .SP4_h_l_00_06(net1377[0:47]),
     .SP12_h_l_00_06(net1378[0:23]), .slf_op_00_06(slf_op_00_06[3:0]),
     .rgt_op_00_06(net1380[0:7]), .SP4_h_l_00_07(net1381[0:47]),
     .SP12_h_l_00_07(net1382[0:23]), .slf_op_00_07(slf_op_00_07[3:0]),
     .rgt_op_00_07(net1384[0:7]), .SP4_h_l_00_08(net1385[0:47]),
     .SP12_h_l_00_08(net1386[0:23]), .slf_op_00_08(slf_op_00_08[3:0]),
     .rgt_op_00_08(slf_op_01_08[7:0]), .fabric_out_01(net1432),
     .fabric_out_02(net1390), .fabric_out_03(net1487),
     .fabric_out_04(net1392), .fabric_out_05(net1478),
     .fabric_out_06(net1479), .fabric_out_07(net1414),
     .fabric_out_08(net1412), .sp4_v_b_00_01(net1397[0:15]),
     .shift(shift_i), .bs_en(bs_en_i), .mode(mode_i), .sdi(sdi),
     .hiz_b(hiz_b_i), .prog(prog), .hold(hold_l_b), .update(update_i),
     .glb_netwk_col(clk_tree_drv[7:0]), .r(r_i), .sdo(net752),
     .bl({bl[0], bl[1], bl[2], bl[3], bl[4], bl[5], bl[6], bl[7],
     bl[8], bl[9], bl[10], bl[11], bl[12], bl[13], bl[14], bl[15],
     bl[16], bl[17]}), .tclk(tclk_i), .ceb(ceb_i));
ice1f_array_BOT_IO_lft12io I_preio_bot_l ( .padin_b_l(padin_b_l[11:0]),
     .padeb_b_l(padeb_b_l[11:0]), .pado_b_l(pado_b_l[11:0]),
     .fabric_out_05_00(net1418), .cf_bot_l(cf_b_l[143:0]),
     .sp4_h_r_06_00(sp4_h_r_06_00[15:0]),
     .tnr_op_06_00(tnr_op_06_00[7:0]), .fabric_out_06_00(net1422),
     .bl_03(bl[167:126]), .bs_en_i(bs_en_bl_1), .ceb_i(ceb_bl_1),
     .hiz_b_i(hiz_b_bl_1), .mode_i(mode_bl_1), .r_i(r_bl_1),
     .shift_i(shift_bl_1), .tclk_i(tclk_bl_1), .update_i(update_bl_1),
     .sdi(sdio_bl_1), .bnl_op_01_00({slf_op_00_01[3], slf_op_00_01[2],
     slf_op_00_01[1], slf_op_00_01[0], slf_op_00_01[3],
     slf_op_00_01[2], slf_op_00_01[1], slf_op_00_01[0]}),
     .sp4_v_b_01_00(net686[0:47]), .slf_op_01_00(slf_op_01_00[3:0]),
     .lft_op_01_00(net1472[0:7]), .sp12_v_b_01_00(net689[0:23]),
     .sp4_v_b_02_00(net690[0:47]), .slf_op_02_00(slf_op_02_00[3:0]),
     .lft_op_02_00(net692[0:7]), .sp12_v_b_02_00(net693[0:23]),
     .sp4_v_b_03_00(net694[0:47]), .slf_op_03_00(slf_op_03_00[3:0]),
     .lft_op_03_00(net696[0:7]), .sp12_v_b_03_00(net697[0:23]),
     .sp4_v_b_04_00(net698[0:47]), .slf_op_04_00(slf_op_04_00[3:0]),
     .lft_op_04_00(net1471[0:7]), .sp12_v_b_04_00(net701[0:23]),
     .sp4_v_b_05_00(net702[0:47]), .slf_op_05_00(slf_op_05_00[3:0]),
     .lft_op_05_00(net704[0:7]), .sp12_v_b_05_00(net705[0:23]),
     .sp4_v_b_06_00(net706[0:47]), .slf_op_06_00(slf_op_06_00[3:0]),
     .lft_op_06_00(slf_op_06_01[7:0]), .sp12_v_b_06_00(net709[0:23]),
     .sp4_h_l_01_00(net1397[0:15]), .hold_b_l(hold_b_l),
     .wl_l({wl_l[1], wl_l[0], wl_l[2], wl_l[3], wl_l[5], wl_l[4],
     wl_l[6], wl_l[7], wl_l[9], wl_l[8], wl_l[10], wl_l[11], wl_l[13],
     wl_l[12], wl_l[14], wl_l[15]}), .vdd_cntl_l({vdd_cntl_l[1],
     vdd_cntl_l[0], vdd_cntl_l[2], vdd_cntl_l[3], vdd_cntl_l[5],
     vdd_cntl_l[4], vdd_cntl_l[6], vdd_cntl_l[7], vdd_cntl_l[9],
     vdd_cntl_l[8], vdd_cntl_l[10], vdd_cntl_l[11], vdd_cntl_l[13],
     vdd_cntl_l[12], vdd_cntl_l[14], vdd_cntl_l[15]}), .tievdd(tievdd),
     .tiegnd(tiegnd), .reset_l({reset_b_l[1], reset_b_l[0],
     reset_b_l[2], reset_b_l[3], reset_b_l[5], reset_b_l[4],
     reset_b_l[6], reset_b_l[7], reset_b_l[9], reset_b_l[8],
     reset_b_l[10], reset_b_l[11], reset_b_l[13], reset_b_l[12],
     reset_b_l[14], reset_b_l[15]}), .prog(prog), .pgate_l({pgate_l[1],
     pgate_l[0], pgate_l[2], pgate_l[3], pgate_l[5], pgate_l[4],
     pgate_l[6], pgate_l[7], pgate_l[9], pgate_l[8], pgate_l[10],
     pgate_l[11], pgate_l[13], pgate_l[12], pgate_l[14], pgate_l[15]}),
     .update_o(update_o), .tclk_o(tclk_o), .shift_o(shift_o),
     .sdo(sdo), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .glb_net_06(net726[0:7]), .glb_net_05(net727[0:7]),
     .glb_net_04(net728[0:7]), .glb_net_03(net729[0:7]),
     .glb_net_02(net730[0:7]), .glb_net_01(net731[0:7]),
     .bs_en_o(bs_en_o), .bl_06(bl[329:276]), .bl_05(bl[275:222]),
     .bl_04(bl[221:168]), .bl_02(bl[125:72]), .bl_01(bl[71:18]),
     .ceb_o(ceb_o));
pinlatbuf12p I_pinlatbuf12p_l ( .pad_in(padin_l_b[13]),
     .icegate(hold_l_b), .cbit(cf_l[183]), .cout(padinlat_l_b[13]),
     .prog(prog));
pinlatbuf12p I_pinlatbuf12p_b ( .pad_in(padin_b_l[11]),
     .icegate(hold_b_l), .cbit(cf_b_l[135]), .cout(padinlat_b_l[11]),
     .prog(prog));
scanbuf1f I_scanbuf_bl ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(net752), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_bl_1), .tclk_o(tclk_bl_1), .shift_o(shift_bl_1),
     .sdo(sdio_bl_1), .r_o(r_bl_1), .mode_o(mode_bl_1),
     .hiz_b_o(hiz_b_bl_1), .ceb_o(ceb_bl_1), .bs_en_o(bs_en_bl_1));
ice1f_array_LT_top I_lt_col_b02 ( .glb_netwk_bo(net730[0:7]),
     .glb_netwk_to(net768[0:7]), .vdd_cntl(vdd_cntl_l[143:16]),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .top_op_08(top_op_02_08[7:0]), .tnl_op_08(tnl_op_02_08[7:0]),
     .tnr_op_08(tnr_op_02_08[7:0]), .sp12_v_t_08(sp12_v_t_02_08[23:0]),
     .sp4_v_t_08(sp4_v_t_02_08[47:0]), .wl(wl_l[143:16]),
     .rgt_op_03(net778[0:7]), .slf_op_02(net1059[0:7]),
     .rgt_op_02(net780[0:7]), .rgt_op_01(net696[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net1372[0:7]), .lft_op_03(net1368[0:7]),
     .lft_op_02(net1364[0:7]), .lft_op_01(net1472[0:7]),
     .rgt_op_04(net788[0:7]), .carry_in(net1486),
     .bnl_op_01({slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0], slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0]}), .slf_op_04(net1067[0:7]),
     .slf_op_03(net1057[0:7]), .slf_op_01(net692[0:7]),
     .sp4_h_l_04(net1086[0:47]), .carry_out(carry_out_02_08),
     .sp12_v_b__01(net693[0:23]), .sp12_h_r_04(net797[0:23]),
     .sp12_h_r_03(net798[0:23]), .sp12_h_r_02(net799[0:23]),
     .sp12_h_r_01(net800[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(net690[0:47]), .sp4_r_v_b_04(net803[0:47]),
     .sp4_r_v_b_03(net804[0:47]), .sp4_r_v_b_02(net805[0:47]),
     .sp4_r_v_b_01(net694[0:47]), .sp4_h_r_04(net807[0:47]),
     .sp4_h_r_03(net808[0:47]), .sp4_h_r_02(net809[0:47]),
     .sp4_h_r_01(net810[0:47]), .sp4_h_l_03(net1087[0:47]),
     .sp4_h_l_02(net1088[0:47]), .sp4_h_l_01(net1089[0:47]),
     .bl(bl[125:72]), .bot_op_01({slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0], slf_op_02_00[3],
     slf_op_02_00[2], slf_op_02_00[1], slf_op_02_00[0]}),
     .sp12_h_l_01(net1079[0:23]), .sp12_h_l_02(net1078[0:23]),
     .sp12_h_l_03(net1077[0:23]), .sp12_h_l_04(net1076[0:23]),
     .sp4_v_b_04(net1082[0:47]), .sp4_v_b_03(net1083[0:47]),
     .sp4_v_b_02(net1084[0:47]), .bnr_op_01({slf_op_03_00[3],
     slf_op_03_00[2], slf_op_03_00[1], slf_op_03_00[0],
     slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0]}), .sp4_h_l_05(net1110[0:47]),
     .sp4_h_l_06(net1109[0:47]), .sp4_h_l_07(net1108[0:47]),
     .sp4_h_l_08(net1107[0:47]), .sp4_h_r_08(net828[0:47]),
     .sp4_h_r_07(net829[0:47]), .sp4_h_r_06(net830[0:47]),
     .sp4_h_r_05(net831[0:47]), .slf_op_05(net1118[0:7]),
     .slf_op_06(net1117[0:7]), .slf_op_07(net1116[0:7]),
     .slf_op_08(slf_op_02_08[7:0]), .rgt_op_08(slf_op_03_08[7:0]),
     .rgt_op_07(net837[0:7]), .rgt_op_06(net838[0:7]),
     .rgt_op_05(net839[0:7]), .lft_op_08(slf_op_01_08[7:0]),
     .lft_op_07(net1384[0:7]), .lft_op_06(net1380[0:7]),
     .lft_op_05(net1376[0:7]), .sp12_h_l_08(net1129[0:23]),
     .sp12_h_l_07(net1128[0:23]), .sp12_h_l_06(net1127[0:23]),
     .sp12_h_r_05(net847[0:23]), .sp12_h_r_06(net848[0:23]),
     .sp12_h_r_07(net849[0:23]), .sp12_h_r_08(net850[0:23]),
     .sp12_h_l_05(net1126[0:23]), .sp4_r_v_b_05(net852[0:47]),
     .sp4_r_v_b_06(net853[0:47]), .sp4_r_v_b_07(net854[0:47]),
     .sp4_r_v_b_08(net855[0:47]), .sp4_v_b_08(net1134[0:47]),
     .sp4_v_b_07(net1133[0:47]), .sp4_v_b_06(net1132[0:47]),
     .sp4_v_b_05(net1131[0:47]));
ice1f_array_LT_top I_lt_col_b06 ( .glb_netwk_bo(net726[0:7]),
     .glb_netwk_to(net1437[0:7]), .vdd_cntl(vdd_cntl_l[143:16]),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .top_op_08(top_op_06_08[7:0]), .tnl_op_08(tnl_op_06_08[7:0]),
     .tnr_op_08(tnr_op_06_08[7:0]), .sp12_v_t_08(sp12_v_t_06_08[23:0]),
     .sp4_v_t_08(sp4_v_t_06_08[47:0]), .wl(wl_l[143:16]),
     .rgt_op_03(rgt_op_06_03[7:0]), .slf_op_02(slf_op_06_02[7:0]),
     .rgt_op_02(rgt_op_06_02[7:0]), .rgt_op_01(rgt_op_06_01[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net974[0:7]),
     .lft_op_03(net964[0:7]), .lft_op_02(net966[0:7]),
     .lft_op_01(net704[0:7]), .rgt_op_04(rgt_op_06_04[7:0]),
     .carry_in(net882), .bnl_op_01({slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0], slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0]}),
     .slf_op_04(slf_op_06_04[7:0]), .slf_op_03(slf_op_06_03[7:0]),
     .slf_op_01(slf_op_06_01[7:0]), .sp4_h_l_04(net1179[0:47]),
     .carry_out(carry_out_06_08), .sp12_v_b__01(net709[0:23]),
     .sp12_h_r_04(sp12_h_r_06_04[23:0]),
     .sp12_h_r_03(sp12_h_r_06_03[23:0]),
     .sp12_h_r_02(sp12_h_r_06_02[23:0]),
     .sp12_h_r_01(sp12_h_r_06_01[23:0]),
     .glb_netwk_col(clk_tree_drv[7:0]), .sp4_v_b_01(net706[0:47]),
     .sp4_r_v_b_04(sp4_r_v_b_06_04[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_06_03[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_06_02[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_06_01[47:0]),
     .sp4_h_r_04(sp4_h_r_06_04[47:0]),
     .sp4_h_r_03(sp4_h_r_06_03[47:0]),
     .sp4_h_r_02(sp4_h_r_06_02[47:0]),
     .sp4_h_r_01(sp4_h_r_06_01[47:0]), .sp4_h_l_03(net1180[0:47]),
     .sp4_h_l_02(net1181[0:47]), .sp4_h_l_01(net1182[0:47]),
     .bl(bl[329:276]), .bot_op_01({slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0], slf_op_06_00[3],
     slf_op_06_00[2], slf_op_06_00[1], slf_op_06_00[0]}),
     .sp12_h_l_01(net1172[0:23]), .sp12_h_l_02(net1171[0:23]),
     .sp12_h_l_03(net1170[0:23]), .sp12_h_l_04(net1169[0:23]),
     .sp4_v_b_04(net1175[0:47]), .sp4_v_b_03(net1176[0:47]),
     .sp4_v_b_02(net1177[0:47]), .bnr_op_01({bnr_op_06_01[3],
     bnr_op_06_01[2], bnr_op_06_01[1], bnr_op_06_01[0],
     bnr_op_06_01[3], bnr_op_06_01[2], bnr_op_06_01[1],
     bnr_op_06_01[0]}), .sp4_h_l_05(net1203[0:47]),
     .sp4_h_l_06(net1202[0:47]), .sp4_h_l_07(net1201[0:47]),
     .sp4_h_l_08(net1200[0:47]), .sp4_h_r_08(sp4_h_r_06_08[47:0]),
     .sp4_h_r_07(sp4_h_r_06_07[47:0]),
     .sp4_h_r_06(sp4_h_r_06_06[47:0]),
     .sp4_h_r_05(sp4_h_r_06_05[47:0]), .slf_op_05(slf_op_06_05[7:0]),
     .slf_op_06(slf_op_06_06[7:0]), .slf_op_07(slf_op_06_07[7:0]),
     .slf_op_08(slf_op_06_08[7:0]), .rgt_op_08(rgt_op_06_08[7:0]),
     .rgt_op_07(rgt_op_06_07[7:0]), .rgt_op_06(rgt_op_06_06[7:0]),
     .rgt_op_05(rgt_op_06_05[7:0]), .lft_op_08(slf_op_05_08[7:0]),
     .lft_op_07(net1023[0:7]), .lft_op_06(net1024[0:7]),
     .lft_op_05(net1025[0:7]), .sp12_h_l_08(net1222[0:23]),
     .sp12_h_l_07(net1221[0:23]), .sp12_h_l_06(net1220[0:23]),
     .sp12_h_r_05(sp12_h_r_06_05[23:0]),
     .sp12_h_r_06(sp12_h_r_06_06[23:0]),
     .sp12_h_r_07(sp12_h_r_06_07[23:0]),
     .sp12_h_r_08(sp12_h_r_06_08[23:0]), .sp12_h_l_05(net1219[0:23]),
     .sp4_r_v_b_05(sp4_r_v_b_06_05[47:0]),
     .sp4_r_v_b_06(sp4_r_v_b_06_06[47:0]),
     .sp4_r_v_b_07(sp4_r_v_b_06_07[47:0]),
     .sp4_r_v_b_08(sp4_r_v_b_06_08[47:0]), .sp4_v_b_08(net1227[0:47]),
     .sp4_v_b_07(net1226[0:47]), .sp4_v_b_06(net1225[0:47]),
     .sp4_v_b_05(net1224[0:47]));
ice1f_array_LT_top I_lt_col_b04 ( .glb_netwk_bo(net728[0:7]),
     .glb_netwk_to(net1452[0:7]), .vdd_cntl(vdd_cntl_l[143:16]),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .top_op_08(top_op_04_08[7:0]), .tnl_op_08(tnl_op_04_08[7:0]),
     .tnr_op_08(tnr_op_04_08[7:0]), .sp12_v_t_08(sp12_v_t_04_08[23:0]),
     .sp4_v_t_08(sp4_v_t_04_08[47:0]), .wl(wl_l[143:16]),
     .rgt_op_03(net964[0:7]), .slf_op_02(net1319[0:7]),
     .rgt_op_02(net966[0:7]), .rgt_op_01(net704[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net788[0:7]), .lft_op_03(net778[0:7]),
     .lft_op_02(net780[0:7]), .lft_op_01(net696[0:7]),
     .rgt_op_04(net974[0:7]), .carry_in(net975),
     .bnl_op_01({slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0], slf_op_03_00[3], slf_op_03_00[2],
     slf_op_03_00[1], slf_op_03_00[0]}), .slf_op_04(net1321[0:7]),
     .slf_op_03(net1318[0:7]), .slf_op_01(net1471[0:7]),
     .sp4_h_l_04(net1330[0:47]), .carry_out(carry_out_04_08),
     .sp12_v_b__01(net701[0:23]), .sp12_h_r_04(net983[0:23]),
     .sp12_h_r_03(net984[0:23]), .sp12_h_r_02(net985[0:23]),
     .sp12_h_r_01(net986[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(net698[0:47]), .sp4_r_v_b_04(net989[0:47]),
     .sp4_r_v_b_03(net990[0:47]), .sp4_r_v_b_02(net991[0:47]),
     .sp4_r_v_b_01(net702[0:47]), .sp4_h_r_04(net993[0:47]),
     .sp4_h_r_03(net994[0:47]), .sp4_h_r_02(net995[0:47]),
     .sp4_h_r_01(net996[0:47]), .sp4_h_l_03(net1331[0:47]),
     .sp4_h_l_02(net1332[0:47]), .sp4_h_l_01(net1333[0:47]),
     .bl(bl[221:168]), .bot_op_01({slf_op_04_00[3], slf_op_04_00[2],
     slf_op_04_00[1], slf_op_04_00[0], slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0]}),
     .sp12_h_l_01(net1305[0:23]), .sp12_h_l_02(net1306[0:23]),
     .sp12_h_l_03(net1267[0:23]), .sp12_h_l_04(net1308[0:23]),
     .sp4_v_b_04(net1283[0:47]), .sp4_v_b_03(net1281[0:47]),
     .sp4_v_b_02(net1279[0:47]), .bnr_op_01({slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0],
     slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0]}), .sp4_h_l_05(net1340[0:47]),
     .sp4_h_l_06(net1338[0:47]), .sp4_h_l_07(net1301[0:47]),
     .sp4_h_l_08(net1302[0:47]), .sp4_h_r_08(net1014[0:47]),
     .sp4_h_r_07(net1015[0:47]), .sp4_h_r_06(net1016[0:47]),
     .sp4_h_r_05(net1017[0:47]), .slf_op_05(net1327[0:7]),
     .slf_op_06(net1328[0:7]), .slf_op_07(net1315[0:7]),
     .slf_op_08(slf_op_04_08[7:0]), .rgt_op_08(slf_op_05_08[7:0]),
     .rgt_op_07(net1023[0:7]), .rgt_op_06(net1024[0:7]),
     .rgt_op_05(net1025[0:7]), .lft_op_08(slf_op_03_08[7:0]),
     .lft_op_07(net837[0:7]), .lft_op_06(net838[0:7]),
     .lft_op_05(net839[0:7]), .sp12_h_l_08(net1266[0:23]),
     .sp12_h_l_07(net1270[0:23]), .sp12_h_l_06(net1263[0:23]),
     .sp12_h_r_05(net1033[0:23]), .sp12_h_r_06(net1034[0:23]),
     .sp12_h_r_07(net1035[0:23]), .sp12_h_r_08(net1036[0:23]),
     .sp12_h_l_05(net1265[0:23]), .sp4_r_v_b_05(net1038[0:47]),
     .sp4_r_v_b_06(net1039[0:47]), .sp4_r_v_b_07(net1040[0:47]),
     .sp4_r_v_b_08(net1041[0:47]), .sp4_v_b_08(net1243[0:47]),
     .sp4_v_b_07(net1303[0:47]), .sp4_v_b_06(net1284[0:47]),
     .sp4_v_b_05(net1286[0:47]));
ice1f_array_LT_top I_lt_col_b01 ( .glb_netwk_bo(net731[0:7]),
     .glb_netwk_to(net1435[0:7]), .vdd_cntl(vdd_cntl_l[143:16]),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .top_op_08(top_op_01_08[7:0]), .tnl_op_08(tnl_op_01_08[7:0]),
     .tnr_op_08(tnr_op_01_08[7:0]), .sp12_v_t_08(sp12_v_t_01_08[23:0]),
     .sp4_v_t_08(sp4_v_t_01_08[47:0]), .wl(wl_l[143:16]),
     .rgt_op_03(net1057[0:7]), .slf_op_02(net1364[0:7]),
     .rgt_op_02(net1059[0:7]), .rgt_op_01(net692[0:7]), .purst(purst),
     .prog(prog), .lft_op_04({slf_op_00_04[3], slf_op_00_04[2],
     slf_op_00_04[1], slf_op_00_04[0], slf_op_00_04[3],
     slf_op_00_04[2], slf_op_00_04[1], slf_op_00_04[0]}),
     .lft_op_03({slf_op_00_03[3], slf_op_00_03[2], slf_op_00_03[1],
     slf_op_00_03[0], slf_op_00_03[3], slf_op_00_03[2],
     slf_op_00_03[1], slf_op_00_03[0]}), .lft_op_02({slf_op_00_02[3],
     slf_op_00_02[2], slf_op_00_02[1], slf_op_00_02[0],
     slf_op_00_02[3], slf_op_00_02[2], slf_op_00_02[1],
     slf_op_00_02[0]}), .lft_op_01({slf_op_00_01[3], slf_op_00_01[2],
     slf_op_00_01[1], slf_op_00_01[0], slf_op_00_01[3],
     slf_op_00_01[2], slf_op_00_01[1], slf_op_00_01[0]}),
     .rgt_op_04(net1067[0:7]), .carry_in(net1068), .bnl_op_01({tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .slf_op_04(net1372[0:7]), .slf_op_03(net1368[0:7]),
     .slf_op_01(net1472[0:7]), .sp4_h_l_04(net1369[0:47]),
     .carry_out(carry_out_01_08), .sp12_v_b__01(net689[0:23]),
     .sp12_h_r_04(net1076[0:23]), .sp12_h_r_03(net1077[0:23]),
     .sp12_h_r_02(net1078[0:23]), .sp12_h_r_01(net1079[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .sp4_v_b_01(net686[0:47]),
     .sp4_r_v_b_04(net1082[0:47]), .sp4_r_v_b_03(net1083[0:47]),
     .sp4_r_v_b_02(net1084[0:47]), .sp4_r_v_b_01(net690[0:47]),
     .sp4_h_r_04(net1086[0:47]), .sp4_h_r_03(net1087[0:47]),
     .sp4_h_r_02(net1088[0:47]), .sp4_h_r_01(net1089[0:47]),
     .sp4_h_l_03(net1365[0:47]), .sp4_h_l_02(net1361[0:47]),
     .sp4_h_l_01(net1466[0:47]), .bl(bl[71:18]),
     .bot_op_01({slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0], slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0]}), .sp12_h_l_01(net1358[0:23]),
     .sp12_h_l_02(net1362[0:23]), .sp12_h_l_03(net1366[0:23]),
     .sp12_h_l_04(net1370[0:23]), .sp4_v_b_04(net1099[0:47]),
     .sp4_v_b_03(net1100[0:47]), .sp4_v_b_02(net1101[0:47]),
     .bnr_op_01({slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0], slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0]}), .sp4_h_l_05(net1373[0:47]),
     .sp4_h_l_06(net1377[0:47]), .sp4_h_l_07(net1381[0:47]),
     .sp4_h_l_08(net1385[0:47]), .sp4_h_r_08(net1107[0:47]),
     .sp4_h_r_07(net1108[0:47]), .sp4_h_r_06(net1109[0:47]),
     .sp4_h_r_05(net1110[0:47]), .slf_op_05(net1376[0:7]),
     .slf_op_06(net1380[0:7]), .slf_op_07(net1384[0:7]),
     .slf_op_08(slf_op_01_08[7:0]), .rgt_op_08(slf_op_02_08[7:0]),
     .rgt_op_07(net1116[0:7]), .rgt_op_06(net1117[0:7]),
     .rgt_op_05(net1118[0:7]), .lft_op_08({slf_op_00_08[3],
     slf_op_00_08[2], slf_op_00_08[1], slf_op_00_08[0],
     slf_op_00_08[3], slf_op_00_08[2], slf_op_00_08[1],
     slf_op_00_08[0]}), .lft_op_07({slf_op_00_07[3], slf_op_00_07[2],
     slf_op_00_07[1], slf_op_00_07[0], slf_op_00_07[3],
     slf_op_00_07[2], slf_op_00_07[1], slf_op_00_07[0]}),
     .lft_op_06({slf_op_00_06[3], slf_op_00_06[2], slf_op_00_06[1],
     slf_op_00_06[0], slf_op_00_06[3], slf_op_00_06[2],
     slf_op_00_06[1], slf_op_00_06[0]}), .lft_op_05({slf_op_00_05[3],
     slf_op_00_05[2], slf_op_00_05[1], slf_op_00_05[0],
     slf_op_00_05[3], slf_op_00_05[2], slf_op_00_05[1],
     slf_op_00_05[0]}), .sp12_h_l_08(net1386[0:23]),
     .sp12_h_l_07(net1382[0:23]), .sp12_h_l_06(net1378[0:23]),
     .sp12_h_r_05(net1126[0:23]), .sp12_h_r_06(net1127[0:23]),
     .sp12_h_r_07(net1128[0:23]), .sp12_h_r_08(net1129[0:23]),
     .sp12_h_l_05(net1374[0:23]), .sp4_r_v_b_05(net1131[0:47]),
     .sp4_r_v_b_06(net1132[0:47]), .sp4_r_v_b_07(net1133[0:47]),
     .sp4_r_v_b_08(net1134[0:47]), .sp4_v_b_08(net1135[0:47]),
     .sp4_v_b_07(net1136[0:47]), .sp4_v_b_06(net1137[0:47]),
     .sp4_v_b_05(net1138[0:47]));
ice1f_array_LT_top I_lt_col_b05 ( .glb_netwk_bo(net727[0:7]),
     .glb_netwk_to(net1453[0:7]), .vdd_cntl(vdd_cntl_l[143:16]),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .top_op_08(top_op_05_08[7:0]), .tnl_op_08(tnl_op_05_08[7:0]),
     .tnr_op_08(tnr_op_05_08[7:0]), .sp12_v_t_08(sp12_v_t_05_08[23:0]),
     .sp4_v_t_08(sp4_v_t_05_08[47:0]), .wl(wl_l[143:16]),
     .rgt_op_03(slf_op_06_03[7:0]), .slf_op_02(net966[0:7]),
     .rgt_op_02(slf_op_06_02[7:0]), .rgt_op_01(slf_op_06_01[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net1321[0:7]),
     .lft_op_03(net1318[0:7]), .lft_op_02(net1319[0:7]),
     .lft_op_01(net1471[0:7]), .rgt_op_04(slf_op_06_04[7:0]),
     .carry_in(net1445), .bnl_op_01({slf_op_04_00[3], slf_op_04_00[2],
     slf_op_04_00[1], slf_op_04_00[0], slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0]}),
     .slf_op_04(net974[0:7]), .slf_op_03(net964[0:7]),
     .slf_op_01(net704[0:7]), .sp4_h_l_04(net993[0:47]),
     .carry_out(carry_out_05_08), .sp12_v_b__01(net705[0:23]),
     .sp12_h_r_04(net1169[0:23]), .sp12_h_r_03(net1170[0:23]),
     .sp12_h_r_02(net1171[0:23]), .sp12_h_r_01(net1172[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .sp4_v_b_01(net702[0:47]),
     .sp4_r_v_b_04(net1175[0:47]), .sp4_r_v_b_03(net1176[0:47]),
     .sp4_r_v_b_02(net1177[0:47]), .sp4_r_v_b_01(net706[0:47]),
     .sp4_h_r_04(net1179[0:47]), .sp4_h_r_03(net1180[0:47]),
     .sp4_h_r_02(net1181[0:47]), .sp4_h_r_01(net1182[0:47]),
     .sp4_h_l_03(net994[0:47]), .sp4_h_l_02(net995[0:47]),
     .sp4_h_l_01(net996[0:47]), .bl(bl[275:222]),
     .bot_op_01({slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0], slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0]}), .sp12_h_l_01(net986[0:23]),
     .sp12_h_l_02(net985[0:23]), .sp12_h_l_03(net984[0:23]),
     .sp12_h_l_04(net983[0:23]), .sp4_v_b_04(net989[0:47]),
     .sp4_v_b_03(net990[0:47]), .sp4_v_b_02(net991[0:47]),
     .bnr_op_01({slf_op_06_00[3], slf_op_06_00[2], slf_op_06_00[1],
     slf_op_06_00[0], slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0]}), .sp4_h_l_05(net1017[0:47]),
     .sp4_h_l_06(net1016[0:47]), .sp4_h_l_07(net1015[0:47]),
     .sp4_h_l_08(net1014[0:47]), .sp4_h_r_08(net1200[0:47]),
     .sp4_h_r_07(net1201[0:47]), .sp4_h_r_06(net1202[0:47]),
     .sp4_h_r_05(net1203[0:47]), .slf_op_05(net1025[0:7]),
     .slf_op_06(net1024[0:7]), .slf_op_07(net1023[0:7]),
     .slf_op_08(slf_op_05_08[7:0]), .rgt_op_08(slf_op_06_08[7:0]),
     .rgt_op_07(slf_op_06_07[7:0]), .rgt_op_06(slf_op_06_06[7:0]),
     .rgt_op_05(slf_op_06_05[7:0]), .lft_op_08(slf_op_04_08[7:0]),
     .lft_op_07(net1315[0:7]), .lft_op_06(net1328[0:7]),
     .lft_op_05(net1327[0:7]), .sp12_h_l_08(net1036[0:23]),
     .sp12_h_l_07(net1035[0:23]), .sp12_h_l_06(net1034[0:23]),
     .sp12_h_r_05(net1219[0:23]), .sp12_h_r_06(net1220[0:23]),
     .sp12_h_r_07(net1221[0:23]), .sp12_h_r_08(net1222[0:23]),
     .sp12_h_l_05(net1033[0:23]), .sp4_r_v_b_05(net1224[0:47]),
     .sp4_r_v_b_06(net1225[0:47]), .sp4_r_v_b_07(net1226[0:47]),
     .sp4_r_v_b_08(net1227[0:47]), .sp4_v_b_08(net1041[0:47]),
     .sp4_v_b_07(net1040[0:47]), .sp4_v_b_06(net1039[0:47]),
     .sp4_v_b_05(net1038[0:47]));
ice1f_array_BRAM_bot I_bram_col_b03 ( .glb_netwk_top(net1428[0:7]),
     .tnr_op_08(tnr_op_03_08[7:0]), .top_op_08(top_op_03_08[7:0]),
     .sp4_v_t_08(sp4_v_t_03_08[47:0]), .tnl_op_08(tnl_op_03_08[7:0]),
     .sp12_v_t_08(sp12_v_t_03_08[23:0]), .pgate(pgate_l[143:16]),
     .reset_b(reset_b_l[143:16]), .vdd_cntl(vdd_cntl_l[143:16]),
     .wl(wl_l[143:16]), .sp4_v_b_08(net855[0:47]),
     .sp4_r_v_b_08(net1243[0:47]), .glb_netwk_bot(net729[0:7]),
     .bm_init_i(bm_init_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sweb_i(bm_sweb_i[1:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sdi_i(bm_sdi_i[1:0]),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sweb_o(bm_sweb_o[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .prog(prog),
     .glb_netwk_col(clk_tree_drv[7:0]), .sp12_h_l_07(net849[0:23]),
     .bnr_op_01({slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0], slf_op_04_00[3], slf_op_04_00[2],
     slf_op_04_00[1], slf_op_04_00[0]}), .sp12_h_r_06(net1263[0:23]),
     .sp12_h_l_06(net848[0:23]), .sp12_h_r_05(net1265[0:23]),
     .sp12_h_r_08(net1266[0:23]), .sp12_h_r_03(net1267[0:23]),
     .sp12_h_l_08(net850[0:23]), .sp12_h_l_05(net847[0:23]),
     .sp12_h_r_07(net1270[0:23]),
     .bm_wdummymux_en_o(bm_wdummymux_en_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .sp4_r_v_b_01(net698[0:47]), .sp4_v_b_02(net805[0:47]),
     .sp4_r_v_b_02(net1279[0:47]), .sp4_v_b_03(net804[0:47]),
     .sp4_r_v_b_03(net1281[0:47]), .sp4_v_b_04(net803[0:47]),
     .sp4_r_v_b_04(net1283[0:47]), .sp4_r_v_b_06(net1284[0:47]),
     .sp4_v_b_06(net853[0:47]), .sp4_r_v_b_05(net1286[0:47]),
     .sp4_v_b_05(net852[0:47]), .lft_op_08(slf_op_02_08[7:0]),
     .lft_op_07(net1116[0:7]), .lft_op_06(net1117[0:7]),
     .lft_op_05(net1118[0:7]), .sp4_v_b_07(net854[0:47]),
     .sp12_h_l_03(net798[0:23]), .sp12_h_l_04(net797[0:23]),
     .sp12_h_l_02(net799[0:23]), .sp12_h_l_01(net800[0:23]),
     .slf_op_07(net837[0:7]), .slf_op_08(slf_op_03_08[7:0]),
     .sp4_h_l_07(net829[0:47]), .sp4_h_l_08(net828[0:47]),
     .sp4_h_r_07(net1301[0:47]), .sp4_h_r_08(net1302[0:47]),
     .sp4_r_v_b_07(net1303[0:47]), .sp4_v_b_01(net694[0:47]),
     .sp12_h_r_01(net1305[0:23]), .sp12_h_r_02(net1306[0:23]),
     .bl(bl[167:126]), .sp12_h_r_04(net1308[0:23]),
     .sp12_v_b_01(net697[0:23]), .bnl_op_01({slf_op_02_00[3],
     slf_op_02_00[2], slf_op_02_00[1], slf_op_02_00[0],
     slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0]}), .lft_op_01(net692[0:7]),
     .lft_op_02(net1059[0:7]), .lft_op_03(net1057[0:7]),
     .lft_op_04(net1067[0:7]), .rgt_op_07(net1315[0:7]),
     .rgt_op_08(slf_op_04_08[7:0]), .bot_op_01({slf_op_03_00[3],
     slf_op_03_00[2], slf_op_03_00[1], slf_op_03_00[0],
     slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0]}), .rgt_op_03(net1318[0:7]),
     .rgt_op_02(net1319[0:7]), .rgt_op_01(net1471[0:7]),
     .rgt_op_04(net1321[0:7]), .slf_op_04(net788[0:7]),
     .slf_op_03(net778[0:7]), .slf_op_02(net780[0:7]),
     .slf_op_01(net696[0:7]), .slf_op_06(net838[0:7]),
     .rgt_op_05(net1327[0:7]), .rgt_op_06(net1328[0:7]),
     .slf_op_05(net839[0:7]), .sp4_h_r_04(net1330[0:47]),
     .sp4_h_r_03(net1331[0:47]), .sp4_h_r_02(net1332[0:47]),
     .sp4_h_r_01(net1333[0:47]), .sp4_h_l_04(net807[0:47]),
     .sp4_h_l_03(net808[0:47]), .sp4_h_l_02(net809[0:47]),
     .sp4_h_l_01(net810[0:47]), .sp4_h_r_06(net1338[0:47]),
     .sp4_h_l_06(net830[0:47]), .sp4_h_r_05(net1340[0:47]),
     .sp4_h_l_05(net831[0:47]));
fabric_outbuf12p I_fbuf_f0008 ( .fabric_out(net1412),
     .cout(fabric_out_00_08));
fabric_outbuf12p I_fbuf_0007 ( .fabric_out(net1414),
     .cout(fabric_out_00_07));
fabric_outbuf12p I_fbuf_p0008b ( .fabric_out(padinlat_l_b[13]),
     .cout(padin_00_08b));
fabric_outbuf12p I_fbuf_f0500 ( .fabric_out(net1418),
     .cout(fabric_out_05_00));
fabric_outbuf12p I_fbuf_p0600b ( .fabric_out(padinlat_b_l[11]),
     .cout(padin_06_00b));
fabric_outbuf12p I_fbuf_f0600 ( .fabric_out(net1422),
     .cout(fabric_out_06_00));
clk_quad_buf12px8 I_clk_quadbuf12px8 ( .clko(clk_tree_drv[7:0]),
     .clki(glb_in[7:0]));

endmodule
// Library - io, Cell - io_col4_RGT_rev, View - schematic
// LAST TIME SAVED: Apr 28 16:05:41 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module io_col4_RGT_rev ( cbit_colcntl, cf, fabric_out, padeb, pado,
     sdo, slf_op, spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l,
     bnl_op, bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op,
     mode, padin, pgate, prog, r, reset, sdi, shift, spioeb, spiout,
     tclk, tnl_op, update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  padeb;
output [23:0]  cf;
output [3:0]  slf_op;
output [1:0]  spi_ss_in_b;
output [1:0]  pado;
output [7:0]  cbit_colcntl;

inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_t;
inout [17:0]  bl;

input [1:0]  spiout;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [7:0]  glb_netwk;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [7:0]  lft_op;
input [15:0]  wl;
input [1:0]  padin;
input [15:0]  reset;
input [1:0]  spioeb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



ioe_col2rev I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .dout(slf_op[3:0]), .outclk(outclk), .hold(hold),
     .rstio(r), .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]}), .reset({reset[14], reset[15], reset[12], reset[13],
     reset[10], reset[11], reset[8], reset[9], reset[6], reset[7],
     reset[4], reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net262), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));
sbox1_colbdlc_rev Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net262));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net262));
rm7  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net262, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .cbit_colcntl(cbit_colcntl[7:0]),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min7({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}), .min5({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14], wl[15],
     wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4],
     wl[5], wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .prog(net262),
     .lc_trk_g1(lc_trk_g1[7:0]));

endmodule
// Library - leafcell, Cell - ice1f_array_RGT_IO_bot9io, View -
//schematic
// LAST TIME SAVED: Aug  3 12:42:33 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module ice1f_array_RGT_IO_bot9io ( cf_r, fabric_out_01, fabric_out_02,
     fabric_out_03, fabric_out_04, fabric_out_05, fabric_out_06,
     fabric_out_07, fabric_out_08, padeb, pado, sdo, slf_op_13_01,
     slf_op_13_02, slf_op_13_03, slf_op_13_04, slf_op_13_05,
     slf_op_13_06, slf_op_13_07, slf_op_13_08, spi_ss_in_b,
     SP4_h_r_13_01, SP4_h_r_13_02, SP4_h_r_13_03, SP4_h_r_13_04,
     SP4_h_r_13_05, SP4_h_r_13_06, SP4_h_r_13_07, SP4_h_r_13_08,
     SP12_h_r_13_01, SP12_h_r_13_02, SP12_h_r_13_03, SP12_h_r_13_04,
     SP12_h_r_13_05, SP12_h_r_13_06, SP12_h_r_13_07, SP12_h_r_13_08,
     bl, pgate, reset_b, sp4_v_b_13_01, sp4_v_t_13_08, vdd_cntl, wl,
     bnl_op_13_01, bs_en, cdone_in, ceb, glb_netwk_col, hiz_b, hold,
     mode, padin, prog, r, rgt_op_13_01, rgt_op_13_02, rgt_op_13_03,
     rgt_op_13_04, rgt_op_13_05, rgt_op_13_06, rgt_op_13_07,
     rgt_op_13_08, sdi, shift, spioeb, spiout, tclk, tnl_op_13_08,
     update );
output  fabric_out_01, fabric_out_02, fabric_out_03, fabric_out_04,
     fabric_out_05, fabric_out_06, fabric_out_07, fabric_out_08, sdo;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_13_01;
output [3:0]  slf_op_13_08;
output [3:0]  slf_op_13_04;
output [3:0]  slf_op_13_02;
output [3:0]  slf_op_13_03;
output [3:0]  slf_op_13_05;
output [15:0]  spi_ss_in_b;
output [8:0]  pado;
output [191:0]  cf_r;
output [3:0]  slf_op_13_06;
output [8:0]  padeb;
output [3:0]  slf_op_13_07;

inout [47:0]  SP4_h_r_13_02;
inout [15:0]  sp4_v_b_13_01;
inout [23:0]  SP12_h_r_13_02;
inout [47:0]  SP4_h_r_13_01;
inout [23:0]  SP12_h_r_13_08;
inout [47:0]  SP4_h_r_13_06;
inout [47:0]  SP4_h_r_13_07;
inout [47:0]  SP4_h_r_13_08;
inout [47:0]  SP4_h_r_13_03;
inout [47:0]  SP4_h_r_13_05;
inout [17:0]  bl;
inout [23:0]  SP12_h_r_13_01;
inout [23:0]  SP12_h_r_13_03;
inout [127:0]  wl;
inout [127:0]  vdd_cntl;
inout [23:0]  SP12_h_r_13_05;
inout [23:0]  SP12_h_r_13_04;
inout [23:0]  SP12_h_r_13_06;
inout [127:0]  pgate;
inout [127:0]  reset_b;
inout [23:0]  SP12_h_r_13_07;
inout [47:0]  SP4_h_r_13_04;
inout [15:0]  sp4_v_t_13_08;

input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_13_01;
input [7:0]  rgt_op_13_04;
input [8:1]  cdone_in;
input [7:0]  tnl_op_13_08;
input [7:0]  rgt_op_13_02;
input [7:0]  rgt_op_13_08;
input [8:0]  padin;
input [15:0]  spioeb;
input [7:0]  rgt_op_13_07;
input [7:0]  rgt_op_13_06;
input [7:0]  rgt_op_13_03;
input [7:0]  rgt_op_13_05;
input [7:0]  bnl_op_13_01;
input [15:0]  spiout;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  noconn00_05;

wire  [0:15]  net486;

wire  [0:15]  net450;

wire  [0:15]  net522;

wire  [0:7]  net635;

wire  [7:0]  glb_netwk_b;

wire  [7:0]  glb_netwk_t;

wire  [7:0]  colbuf_cntl_b;

wire  [7:0]  colbuf_cntl_t;

wire  [0:15]  net414;

wire  [0:1]  net520;

wire  [0:15]  net594;

wire  [0:1]  net485;

wire  [0:7]  net636;

wire  [0:1]  net521;

wire  [0:7]  net628;

wire  [0:7]  net638;

wire  [0:15]  net378;

wire  [0:7]  net541;

wire  [0:1]  net484;

wire  [0:1]  net0623;

wire  [0:7]  net629;

wire  [0:15]  net558;



io_col4_RGT_rev I_io_00_08 ( .cbit_colcntl(net629[0:7]), .ceb(ceb),
     .sdo(sdo), .sdi(net363), .spiout(spiout[15:14]),
     .cdone_in(cdone_in[8]), .spioeb(spioeb[15:14]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[8:7]), .pado(pado[8:7]),
     .padeb(padeb[8:7]), .sp4_v_t(sp4_v_t_13_08[15:0]),
     .sp4_h_l(SP4_h_r_13_08[47:0]), .sp12_h_l(SP12_h_r_13_08[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[15:14]),
     .tnl_op(tnl_op_13_08[7:0]), .lft_op(rgt_op_13_08[7:0]),
     .bnl_op(rgt_op_13_07[7:0]), .pgate(pgate[127:112]),
     .reset(reset_b[127:112]), .sp4_v_b(net378[0:15]),
     .wl(wl[127:112]), .cf(cf_r[191:168]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[127:112]), .slf_op(slf_op_13_08[3:0]),
     .glb_netwk(glb_netwk_t[7:0]), .hold(hold),
     .fabric_out(fabric_out_08));
io_col4_RGT_rev I_io_00_07 ( .cbit_colcntl(net636[0:7]), .ceb(ceb),
     .sdo(net363), .sdi(net435), .spiout(spiout[13:12]),
     .cdone_in(cdone_in[7]), .spioeb(spioeb[13:12]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[6:5]), .pado(pado[6:5]),
     .padeb(padeb[6:5]), .sp4_v_t(net378[0:15]),
     .sp4_h_l(SP4_h_r_13_07[47:0]), .sp12_h_l(SP12_h_r_13_07[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[13:12]),
     .tnl_op(rgt_op_13_08[7:0]), .lft_op(rgt_op_13_07[7:0]),
     .bnl_op(rgt_op_13_06[7:0]), .pgate(pgate[111:96]),
     .reset(reset_b[111:96]), .sp4_v_b(net450[0:15]), .wl(wl[111:96]),
     .cf(cf_r[167:144]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_13_07[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_07));
io_col4_RGT_rev I_io_00_05 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net399), .sdi(net579), .spiout(spiout[9:8]),
     .cdone_in(cdone_in[5]), .spioeb(spioeb[9:8]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(noconn00_05[1:0]),
     .pado(noconn00_05[1:0]), .padeb(net0623[0:1]),
     .sp4_v_t(net414[0:15]), .sp4_h_l(SP4_h_r_13_05[47:0]),
     .sp12_h_l(SP12_h_r_13_05[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[9:8]), .tnl_op(rgt_op_13_06[7:0]),
     .lft_op(rgt_op_13_05[7:0]), .bnl_op(rgt_op_13_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net594[0:15]), .wl(wl[79:64]), .cf(cf_r[119:96]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_13_05[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_05));
io_col4_RGT_rev I_io_00_06 ( .cbit_colcntl(net638[0:7]), .ceb(ceb),
     .sdo(net435), .sdi(net399), .spiout(spiout[11:10]),
     .cdone_in(cdone_in[6]), .spioeb(spioeb[11:10]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[4:3]), .pado(pado[4:3]),
     .padeb(padeb[4:3]), .sp4_v_t(net450[0:15]),
     .sp4_h_l(SP4_h_r_13_06[47:0]), .sp12_h_l(SP12_h_r_13_06[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[11:10]),
     .tnl_op(rgt_op_13_07[7:0]), .lft_op(rgt_op_13_06[7:0]),
     .bnl_op(rgt_op_13_05[7:0]), .pgate(pgate[95:80]),
     .reset(reset_b[95:80]), .sp4_v_b(net414[0:15]), .wl(wl[95:80]),
     .cf(cf_r[143:120]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_13_06[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_06));
io_col4_RGT_rev I_io_00_02 ( .cbit_colcntl(net628[0:7]), .ceb(ceb),
     .sdo(net471), .sdi(net507), .spiout(spiout[3:2]),
     .cdone_in(cdone_in[2]), .spioeb(spioeb[3:2]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(net484[0:1]), .pado(net484[0:1]),
     .padeb(net485[0:1]), .sp4_v_t(net486[0:15]),
     .sp4_h_l(SP4_h_r_13_02[47:0]), .sp12_h_l(SP12_h_r_13_02[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[3:2]),
     .tnl_op(rgt_op_13_03[7:0]), .lft_op(rgt_op_13_02[7:0]),
     .bnl_op(rgt_op_13_01[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b(net522[0:15]), .wl(wl[31:16]),
     .cf(cf_r[47:24]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_13_02[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_02));
io_col4_RGT_rev I_io_00_01 ( .cbit_colcntl(net635[0:7]), .ceb(ceb),
     .sdo(net507), .sdi(sdi), .spiout(spiout[1:0]),
     .cdone_in(cdone_in[1]), .spioeb(spioeb[1:0]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(net520[0:1]), .pado(net520[0:1]),
     .padeb(net521[0:1]), .sp4_v_t(net522[0:15]),
     .sp4_h_l(SP4_h_r_13_01[47:0]), .sp12_h_l(SP12_h_r_13_01[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[1:0]),
     .tnl_op(rgt_op_13_02[7:0]), .lft_op(rgt_op_13_01[7:0]),
     .bnl_op(bnl_op_13_01[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(sp4_v_b_13_01[15:0]),
     .wl(wl[15:0]), .cf(cf_r[23:0]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_13_01[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold),
     .fabric_out(fabric_out_01));
io_col4_RGT_rev I_io_00_03 ( .cbit_colcntl(net541[0:7]), .ceb(ceb),
     .sdo(net543), .sdi(net471), .spiout(spiout[5:4]),
     .cdone_in(cdone_in[3]), .spioeb(spioeb[5:4]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin({padin[0], padin0off}), .pado({pado[0],
     padin0off}), .padeb({padeb[0], padeb0off}),
     .sp4_v_t(net558[0:15]), .sp4_h_l(SP4_h_r_13_03[47:0]),
     .sp12_h_l(SP12_h_r_13_03[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[5:4]), .tnl_op(rgt_op_13_04[7:0]),
     .lft_op(rgt_op_13_03[7:0]), .bnl_op(rgt_op_13_02[7:0]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net486[0:15]), .wl(wl[47:32]), .cf(cf_r[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_13_03[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_03));
io_col4_RGT_rev I_io_00_04 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net579), .sdi(net543), .spiout(spiout[7:6]),
     .cdone_in(cdone_in[4]), .spioeb(spioeb[7:6]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[2:1]), .pado(pado[2:1]),
     .padeb(padeb[2:1]), .sp4_v_t(net594[0:15]),
     .sp4_h_l(SP4_h_r_13_04[47:0]), .sp12_h_l(SP12_h_r_13_04[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[7:6]),
     .tnl_op(rgt_op_13_05[7:0]), .lft_op(rgt_op_13_04[7:0]),
     .bnl_op(rgt_op_13_03[7:0]), .pgate(pgate[63:48]),
     .reset(reset_b[63:48]), .sp4_v_b(net558[0:15]), .wl(wl[63:48]),
     .cf(cf_r[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_13_04[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_04));
clk_colbuf1kx8 Iclk_colbuf1kx8_t ( .colbuf_cntl(colbuf_cntl_t[7:0]),
     .col_clk(glb_netwk_t[7:0]), .clk_in(glb_netwk_col[7:0]));
clk_colbuf1kx8 I_clk_colbuf1kx8_b ( .colbuf_cntl(colbuf_cntl_b[7:0]),
     .col_clk(glb_netwk_b[7:0]), .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - leafcell, Cell - ice1f_array_BOT_IO_rgt12io, View -
//schematic
// LAST TIME SAVED: Jul 16 17:13:07 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module ice1f_array_BOT_IO_rgt12io ( cf_bot_r, fabric_out_07_00,
     fabric_out_12_00, padeb_b_r, pado_b_r, sdo, slf_op_01_00,
     slf_op_02_00, slf_op_03_00, slf_op_04_00, slf_op_05_00,
     slf_op_06_00, spi_ss_in_b, bl_01, bl_02, bl_03, bl_04, bl_05,
     bl_06, sp4_h_l_21_00, sp4_h_r_06_00, sp4_v_b_01_00, sp4_v_b_02_00,
     sp4_v_b_03_00, sp4_v_b_04_00, sp4_v_b_05_00, sp4_v_b_06_00,
     sp12_v_b_01_00, sp12_v_b_02_00, sp12_v_b_03_00, sp12_v_b_04_00,
     sp12_v_b_05_00, sp12_v_b_06_00, bnl_op_01_00, bs_en_i, ceb_i,
     end_of_startup_top_l, glb_net_01, glb_net_02, glb_net_03,
     glb_net_04, glb_net_05, glb_net_06, hiz_b_i, hold_b_r,
     lft_op_01_00, lft_op_02_00, lft_op_03_00, lft_op_04_00,
     lft_op_05_00, lft_op_06_00, mode_i, padin_b_r, pgate_l, prog, r_i,
     reset_l, sdi, shift_i, spiceb, spiout, tclk_i, tnr_op_06_00,
     update_i, vdd_cntl_l, wl_l );
output  fabric_out_07_00, fabric_out_12_00, sdo;


input  bs_en_i, ceb_i, hiz_b_i, hold_b_r, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_05_00;
output [11:0]  spi_ss_in_b;
output [143:0]  cf_bot_r;
output [11:0]  padeb_b_r;
output [11:0]  pado_b_r;
output [3:0]  slf_op_04_00;
output [3:0]  slf_op_02_00;
output [3:0]  slf_op_01_00;
output [3:0]  slf_op_03_00;
output [3:0]  slf_op_06_00;

inout [47:0]  sp4_v_b_01_00;
inout [47:0]  sp4_v_b_02_00;
inout [23:0]  sp12_v_b_05_00;
inout [47:0]  sp4_v_b_03_00;
inout [23:0]  sp12_v_b_03_00;
inout [47:0]  sp4_v_b_04_00;
inout [23:0]  sp12_v_b_01_00;
inout [23:0]  sp12_v_b_04_00;
inout [23:0]  sp12_v_b_06_00;
inout [41:0]  bl_04;
inout [53:0]  bl_05;
inout [53:0]  bl_02;
inout [53:0]  bl_03;
inout [53:0]  bl_01;
inout [15:0]  sp4_h_l_21_00;
inout [23:0]  sp12_v_b_02_00;
inout [47:0]  sp4_v_b_06_00;
inout [15:0]  sp4_h_r_06_00;
inout [53:0]  bl_06;
inout [47:0]  sp4_v_b_05_00;

input [7:0]  glb_net_03;
input [7:0]  glb_net_05;
input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_01;
input [7:0]  bnl_op_01_00;
input [7:0]  tnr_op_06_00;
input [7:0]  lft_op_04_00;
input [7:0]  lft_op_06_00;
input [15:0]  pgate_l;
input [7:0]  lft_op_02_00;
input [11:0]  spiceb;
input [11:0]  spiout;
input [6:1]  end_of_startup_top_l;
input [11:0]  padin_b_r;
input [15:0]  wl_l;
input [7:0]  glb_net_06;
input [7:0]  lft_op_01_00;
input [7:0]  lft_op_03_00;
input [15:0]  reset_l;
input [7:0]  lft_op_05_00;
input [7:0]  glb_net_02;
input [7:0]  glb_net_04;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net379;

wire  [0:15]  net309;

wire  [0:15]  net414;

wire  [0:15]  net344;

wire  [0:15]  net274;



io_col4_BOT_rev I_io_b07 ( .sdo(net258), .sdi(sdi),
     .spiout(spiout[1:0]), .cdone_in(end_of_startup_top_l[1]),
     .spioeb(spiceb[1:0]), .sp4_v_t(sp4_h_l_21_00[15:0]),
     .mode(mode_i), .shift(shift_i), .hiz_b(hiz_b_i), .r(r_i),
     .bs_en(bs_en_i), .tclk(tclk_i), .update(update_i),
     .padin(padin_b_r[1:0]), .pado(pado_b_r[1:0]),
     .padeb(padeb_b_r[1:0]), .sp4_v_b(net274[0:15]),
     .sp4_h_l(sp4_v_b_01_00[47:0]), .sp12_h_l(sp12_v_b_01_00[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[1:0]),
     .tnl_op(bnl_op_01_00[7:0]), .lft_op(lft_op_01_00[7:0]),
     .bnl_op(lft_op_02_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_r[23:0]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_00[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_b_r), .fabric_out(fabric_out_07_00));
io_col4_BOT_rev I_io_b08 ( .sdo(net293), .sdi(net258),
     .spiout(spiout[3:2]), .cdone_in(end_of_startup_top_l[2]),
     .spioeb(spiceb[3:2]), .sp4_v_t(net274[0:15]), .mode(mode_i),
     .shift(shift_i), .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i),
     .tclk(tclk_i), .update(update_i), .padin(padin_b_r[3:2]),
     .pado(pado_b_r[3:2]), .padeb(padeb_b_r[3:2]),
     .sp4_v_b(net309[0:15]), .sp4_h_l(sp4_v_b_02_00[47:0]),
     .sp12_h_l(sp12_v_b_02_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[3:2]), .tnl_op(lft_op_01_00[7:0]),
     .lft_op(lft_op_02_00[7:0]), .bnl_op(lft_op_03_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_02[5],
     bl_02[4], bl_02[37], bl_02[36], bl_02[35], bl_02[34], bl_02[33],
     bl_02[32], bl_02[14], bl_02[20], bl_02[19], bl_02[18], bl_02[17],
     bl_02[16], bl_02[27], bl_02[26], bl_02[25], bl_02[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_r[47:24]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_02_00[3:0]),
     .glb_netwk(glb_net_02[7:0]), .hold(hold_b_r),
     .fabric_out(net327));
io_col4_BOT_rev I_io_b09 ( .sdo(net328), .sdi(net293),
     .spiout(spiout[5:4]), .cdone_in(end_of_startup_top_l[3]),
     .spioeb(spiceb[5:4]), .sp4_v_t(net309[0:15]), .mode(mode_i),
     .shift(shift_i), .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i),
     .tclk(tclk_i), .update(update_i), .padin(padin_b_r[5:4]),
     .pado(pado_b_r[5:4]), .padeb(padeb_b_r[5:4]),
     .sp4_v_b(net344[0:15]), .sp4_h_l(sp4_v_b_03_00[47:0]),
     .sp12_h_l(sp12_v_b_03_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[5:4]), .tnl_op(lft_op_02_00[7:0]),
     .lft_op(lft_op_03_00[7:0]), .bnl_op(lft_op_04_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_03[5],
     bl_03[4], bl_03[37], bl_03[36], bl_03[35], bl_03[34], bl_03[33],
     bl_03[32], bl_03[14], bl_03[20], bl_03[19], bl_03[18], bl_03[17],
     bl_03[16], bl_03[27], bl_03[26], bl_03[25], bl_03[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_r[71:48]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_03_00[3:0]),
     .glb_netwk(glb_net_03[7:0]), .hold(hold_b_r),
     .fabric_out(net362));
io_col4_BOT_rev I_io_b11 ( .sdo(net363), .sdi(net398),
     .spiout(spiout[9:8]), .cdone_in(end_of_startup_top_l[5]),
     .spioeb(spiceb[9:8]), .sp4_v_t(net414[0:15]), .mode(mode_i),
     .shift(shift_i), .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i),
     .tclk(tclk_i), .update(update_i), .padin(padin_b_r[9:8]),
     .pado(pado_b_r[9:8]), .padeb(padeb_b_r[9:8]),
     .sp4_v_b(net379[0:15]), .sp4_h_l(sp4_v_b_05_00[47:0]),
     .sp12_h_l(sp12_v_b_05_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[9:8]), .tnl_op(lft_op_04_00[7:0]),
     .lft_op(lft_op_05_00[7:0]), .bnl_op(lft_op_06_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_05[5],
     bl_05[4], bl_05[37], bl_05[36], bl_05[35], bl_05[34], bl_05[33],
     bl_05[32], bl_05[14], bl_05[20], bl_05[19], bl_05[18], bl_05[17],
     bl_05[16], bl_05[27], bl_05[26], bl_05[25], bl_05[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_r[119:96]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_05_00[3:0]),
     .glb_netwk(glb_net_05[7:0]), .hold(hold_b_r),
     .fabric_out(net483));
io_col4_BOT_rev I_io_b10 ( .sdo(net398), .sdi(net328),
     .spiout(spiout[7:6]), .cdone_in(end_of_startup_top_l[4]),
     .spioeb(spiceb[7:6]), .sp4_v_t(net344[0:15]), .mode(mode_i),
     .shift(shift_i), .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i),
     .tclk(tclk_i), .update(update_i), .padin(padin_b_r[7:6]),
     .pado(pado_b_r[7:6]), .padeb(padeb_b_r[7:6]),
     .sp4_v_b(net414[0:15]), .sp4_h_l(sp4_v_b_04_00[47:0]),
     .sp12_h_l(sp12_v_b_04_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[7:6]), .tnl_op(lft_op_03_00[7:0]),
     .lft_op(lft_op_04_00[7:0]), .bnl_op(lft_op_05_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_04[5],
     bl_04[4], bl_04[37], bl_04[36], bl_04[35], bl_04[34], bl_04[33],
     bl_04[32], bl_04[14], bl_04[20], bl_04[19], bl_04[18], bl_04[17],
     bl_04[16], bl_04[27], bl_04[26], bl_04[25], bl_04[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_r[95:72]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_04_00[3:0]),
     .glb_netwk(glb_net_04[7:0]), .hold(hold_b_r),
     .fabric_out(net432));
io_col4_BOT_rev I_io_b12 ( .sdo(net433), .sdi(net363),
     .spiout(spiout[11:10]), .cdone_in(end_of_startup_top_l[6]),
     .spioeb(spiceb[11:10]), .sp4_v_t(net379[0:15]), .mode(mode_i),
     .shift(shift_i), .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i),
     .tclk(tclk_i), .update(update_i), .padin(padin_b_r[11:10]),
     .pado(pado_b_r[11:10]), .padeb(padeb_b_r[11:10]),
     .sp4_v_b(sp4_h_r_06_00[15:0]), .sp4_h_l(sp4_v_b_06_00[47:0]),
     .sp12_h_l(sp12_v_b_06_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[11:10]), .tnl_op(lft_op_05_00[7:0]),
     .lft_op(lft_op_06_00[7:0]), .bnl_op(tnr_op_06_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_06[5],
     bl_06[4], bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33],
     bl_06[32], bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17],
     bl_06[16], bl_06[27], bl_06[26], bl_06[25], bl_06[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_r[143:120]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_06_00[3:0]),
     .glb_netwk(glb_net_06[7:0]), .hold(hold_b_r),
     .fabric_out(fabric_out_12_00));
lowla_modified I_lowla_brout ( .clk(tclk_i), .min(net257), .lao(sdo));
bram_bufferx4x6 I_sdibuf ( .in(net433), .out(net257));

endmodule
// Library - leafcell, Cell - ice1f_quad_br, View - schematic
// LAST TIME SAVED: Jul 22 09:50:59 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module ice1f_quad_br ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_07_08, carry_out_08_08,
     carry_out_09_08, carry_out_11_08, carry_out_12_08, ceb_o, cf_b,
     cf_r, fabric_out_07_00, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fabric_out_13_08, hiz_b_o, mode_o, padeb_b_r,
     padeb_r_b, padin_07_00a, padin_13_08b, pado_b_r, pado_r_b, r_o,
     sdo, sdo_pad, shift_o, slf_op_07_00, slf_op_07_01, slf_op_07_02,
     slf_op_07_03, slf_op_07_04, slf_op_07_05, slf_op_07_06,
     slf_op_07_07, slf_op_07_08, slf_op_08_08, slf_op_09_08,
     slf_op_10_08, slf_op_11_08, slf_op_12_08, slf_op_13_08,
     spi_ss_in_b, spi_ss_in_r, tclk_o, update_o, bl, pgate_r,
     reset_b_r, sp4_h_l_07_00, sp4_h_l_07_01, sp4_h_l_07_02,
     sp4_h_l_07_03, sp4_h_l_07_04, sp4_h_l_07_05, sp4_h_l_07_06,
     sp4_h_l_07_07, sp4_h_l_07_08, sp4_v_b_07_01, sp4_v_b_07_02,
     sp4_v_b_07_03, sp4_v_b_07_04, sp4_v_b_07_05, sp4_v_b_07_06,
     sp4_v_b_07_07, sp4_v_b_07_08, sp4_v_t_07_08, sp4_v_t_08_08,
     sp4_v_t_09_08, sp4_v_t_10_08, sp4_v_t_11_08, sp4_v_t_12_08,
     sp4_v_t_13_08, sp12_h_l_07_01, sp12_h_l_07_02, sp12_h_l_07_03,
     sp12_h_l_07_04, sp12_h_l_07_05, sp12_h_l_07_06, sp12_h_l_07_07,
     sp12_h_l_07_08, sp12_v_t_07_08, sp12_v_t_08_08, sp12_v_t_09_08,
     sp12_v_t_10_08, sp12_v_t_11_08, sp12_v_t_12_08, vdd_cntl_r, wl_r,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i,
     bnl_op_07_01, bs_en_i, bs_en_mi, ceb_i, ceb_mi,
     end_of_startup_bot_r, end_of_startup_rgt_b, glb_in, hiz_b_i,
     hiz_b_mi, hold_b_r, hold_r_b, mode_i, mode_mi, padin_b_r,
     padin_r_b, prog, purst, r_i, r_mi, rgt_op_07_01, rgt_op_07_02,
     rgt_op_07_03, rgt_op_07_04, rgt_op_07_05, rgt_op_07_06,
     rgt_op_07_07, rgt_op_07_08, sdi, sdi_pad, shift_i, shift_mi,
     spioeb, spioeb_r, spiout, spiout_r, tclk_i, tclk_mi, tiegnd,
     tnl_op_07_08, tnl_op_08_08, tnl_op_09_08, tnl_op_10_08,
     tnl_op_11_08, tnl_op_12_08, tnr_op_07_08, tnr_op_08_08,
     tnr_op_09_08, tnr_op_10_08, tnr_op_11_08, tnr_op_12_08,
     top_op_07_08, top_op_08_08, top_op_09_08, top_op_10_08,
     top_op_11_08, top_op_12_08, update_i, update_mi );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_07_08, carry_out_08_08,
     carry_out_09_08, carry_out_11_08, carry_out_12_08, ceb_o,
     fabric_out_07_00, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fabric_out_13_08, hiz_b_o, mode_o, padin_07_00a,
     padin_13_08b, r_o, sdo, sdo_pad, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, bs_en_mi, ceb_i, ceb_mi, hiz_b_i,
     hiz_b_mi, hold_b_r, hold_r_b, mode_i, mode_mi, prog, purst, r_i,
     r_mi, sdi, sdi_pad, shift_i, shift_mi, tclk_i, tclk_mi, tiegnd,
     update_i, update_mi;

output [1:0]  bm_sweb_o;
output [7:0]  slf_op_08_08;
output [7:0]  slf_op_07_02;
output [3:0]  slf_op_07_00;
output [8:0]  pado_r_b;
output [8:0]  padeb_r_b;
output [15:0]  spi_ss_in_r;
output [11:0]  padeb_b_r;
output [7:0]  slf_op_11_08;
output [7:0]  slf_op_07_07;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_07_04;
output [7:0]  slf_op_10_08;
output [3:0]  slf_op_13_08;
output [7:0]  slf_op_07_05;
output [7:0]  slf_op_07_06;
output [11:0]  pado_b_r;
output [1:0]  bm_sdo_o;
output [11:0]  spi_ss_in_b;
output [1:0]  bm_sdi_o;
output [143:0]  cf_b;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_07_01;
output [7:0]  slf_op_07_03;
output [7:0]  slf_op_07_08;
output [7:0]  slf_op_12_08;
output [191:0]  cf_r;
output [7:0]  slf_op_09_08;

inout [47:0]  sp4_v_t_09_08;
inout [47:0]  sp4_h_l_07_01;
inout [47:0]  sp4_h_l_07_04;
inout [23:0]  sp12_h_l_07_06;
inout [47:0]  sp4_v_t_12_08;
inout [23:0]  sp12_h_l_07_03;
inout [47:0]  sp4_h_l_07_05;
inout [47:0]  sp4_v_t_08_08;
inout [47:0]  sp4_v_t_10_08;
inout [47:0]  sp4_h_l_07_06;
inout [47:0]  sp4_v_t_11_08;
inout [23:0]  sp12_h_l_07_02;
inout [47:0]  sp4_v_b_07_02;
inout [23:0]  sp12_h_l_07_07;
inout [23:0]  sp12_v_t_07_08;
inout [143:0]  pgate_r;
inout [23:0]  sp12_v_t_10_08;
inout [23:0]  sp12_v_t_08_08;
inout [23:0]  sp12_v_t_11_08;
inout [47:0]  sp4_v_b_07_07;
inout [47:0]  sp4_v_b_07_03;
inout [47:0]  sp4_v_b_07_08;
inout [47:0]  sp4_h_l_07_07;
inout [47:0]  sp4_h_l_07_02;
inout [47:0]  sp4_v_b_07_06;
inout [47:0]  sp4_v_b_07_05;
inout [23:0]  sp12_v_t_12_08;
inout [23:0]  sp12_h_l_07_08;
inout [47:0]  sp4_v_b_07_01;
inout [143:0]  wl_r;
inout [23:0]  sp12_h_l_07_04;
inout [47:0]  sp4_h_l_07_08;
inout [47:0]  sp4_h_l_07_03;
inout [47:0]  sp4_v_b_07_04;
inout [47:0]  sp4_v_t_07_08;
inout [329:0]  bl;
inout [15:0]  sp4_h_l_07_00;
inout [143:0]  reset_b_r;
inout [15:0]  sp4_v_t_13_08;
inout [143:0]  vdd_cntl_r;
inout [23:0]  sp12_v_t_09_08;
inout [23:0]  sp12_h_l_07_05;
inout [23:0]  sp12_h_l_07_01;

input [7:0]  top_op_09_08;
input [7:0]  rgt_op_07_02;
input [7:0]  top_op_12_08;
input [7:0]  top_op_08_08;
input [7:0]  rgt_op_07_03;
input [7:0]  bm_sa_i;
input [7:0]  rgt_op_07_08;
input [15:0]  spioeb_r;
input [11:0]  spioeb;
input [7:0]  tnl_op_09_08;
input [7:0]  tnl_op_11_08;
input [7:0]  tnr_op_12_08;
input [7:0]  tnl_op_10_08;
input [7:0]  tnl_op_07_08;
input [7:0]  top_op_11_08;
input [7:0]  rgt_op_07_05;
input [7:0]  rgt_op_07_07;
input [7:0]  rgt_op_07_06;
input [7:0]  rgt_op_07_04;
input [1:0]  bm_sclkrw_i;
input [15:0]  spiout_r;
input [7:0]  glb_in;
input [7:0]  tnl_op_12_08;
input [7:0]  rgt_op_07_01;
input [7:0]  tnr_op_11_08;
input [11:0]  spiout;
input [7:0]  tnr_op_07_08;
input [7:0]  tnr_op_10_08;
input [1:0]  bm_sweb_i;
input [8:0]  padin_r_b;
input [3:0]  bnl_op_07_01;
input [7:0]  tnr_op_09_08;
input [1:0]  bm_sdi_i;
input [11:0]  padin_b_r;
input [8:1]  end_of_startup_rgt_b;
input [7:0]  top_op_10_08;
input [7:0]  tnl_op_08_08;
input [7:0]  top_op_07_08;
input [1:0]  bm_sdo_i;
input [7:0]  tnr_op_08_08;
input [12:7]  end_of_startup_bot_r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net1049;

wire  [0:47]  net834;

wire  [0:47]  net1225;

wire  [0:7]  net0855;

wire  [0:47]  net1385;

wire  [0:47]  net1382;

wire  [0:47]  net969;

wire  [0:47]  net1294;

wire  [0:23]  net1377;

wire  [0:7]  net1142;

wire  [0:7]  net1233;

wire  [0:7]  net858;

wire  [0:7]  net1493;

wire  [0:7]  net0859;

wire  [0:47]  net1290;

wire  [0:7]  net1081;

wire  [0:23]  net1284;

wire  [0:7]  net862;

wire  [0:47]  net1132;

wire  [0:7]  net828;

wire  [0:47]  net1340;

wire  [0:47]  net978;

wire  [0:47]  net1108;

wire  [0:7]  net1048;

wire  [7:0]  clk_tree_drv;

wire  [0:47]  net1014;

wire  [0:47]  net939;

wire  [0:7]  net965;

wire  [0:15]  net811;

wire  [0:23]  net1152;

wire  [0:7]  net1050;

wire  [0:23]  net1195;

wire  [0:23]  net904;

wire  [0:7]  net957;

wire  [3:0]  slf_op_12_00;

wire  [0:47]  net938;

wire  [0:47]  net971;

wire  [0:23]  net1334;

wire  [0:23]  net1150;

wire  [0:47]  net1064;

wire  [0:47]  net918;

wire  [0:47]  net1291;

wire  [0:7]  net1326;

wire  [0:47]  net1480;

wire  [0:47]  net1200;

wire  [0:23]  net1376;

wire  [0:7]  net989;

wire  [0:7]  net1083;

wire  [0:23]  net837;

wire  [0:23]  net1151;

wire  [0:47]  net1317;

wire  [0:47]  net968;

wire  [0:47]  net1112;

wire  [0:47]  net1250;

wire  [0:23]  net1287;

wire  [0:47]  net1107;

wire  [0:23]  net833;

wire  [0:7]  net1091;

wire  [0:47]  net1297;

wire  [0:47]  net1481;

wire  [0:47]  net941;

wire  [0:23]  net1245;

wire  [11:11]  padinlat_r_b;

wire  [0:23]  net1285;

wire  [0:47]  net1496;

wire  [0:7]  net0860;

wire  [0:7]  net863;

wire  [0:47]  net1134;

wire  [0:47]  net1384;

wire  [0:47]  net1016;

wire  [0:23]  net1100;

wire  [0:7]  net1140;

wire  [0:47]  net1223;

wire  [0:47]  net1339;

wire  [0:23]  net1193;

wire  [0:23]  net1060;

wire  [0:23]  net1058;

wire  [0:47]  net1113;

wire  [0:47]  net1248;

wire  [0:23]  net1244;

wire  [0:47]  net1110;

wire  [0:7]  net1141;

wire  [0:23]  net1426;

wire  [0:23]  net1286;

wire  [0:23]  net1428;

wire  [0:7]  net859;

wire  [3:0]  slf_op_13_07;

wire  [0:23]  net907;

wire  [0:7]  net836;

wire  [0:47]  net1199;

wire  [0:23]  net903;

wire  [0:47]  net1431;

wire  [0:47]  net1155;

wire  [0:23]  net1009;

wire  [0:23]  net1242;

wire  [0:47]  net1224;

wire  [0:7]  net0856;

wire  [0:47]  net1204;

wire  [0:47]  net1156;

wire  [0:47]  net1433;

wire  [0:47]  net970;

wire  [0:23]  net1194;

wire  [0:47]  net1202;

wire  [0:47]  net1018;

wire  [0:47]  net1434;

wire  [0:47]  net1131;

wire  [0:47]  net1506;

wire  [0:47]  net1407;

wire  [0:23]  net1192;

wire  [0:23]  net944;

wire  [0:47]  net1040;

wire  [0:7]  net1267;

wire  [0:7]  net1232;

wire  [0:47]  net1318;

wire  [0:47]  net976;

wire  [0:47]  net1342;

wire  [0:23]  net1379;

wire  [0:7]  net1275;

wire  [0:47]  net1063;

wire  [0:47]  net1041;

wire  [0:47]  net1295;

wire  [0:7]  net1175;

wire  [3:0]  slf_op_13_02;

wire  [3:0]  slf_op_13_01;

wire  [0:47]  net1383;

wire  [0:23]  net1243;

wire  [0:23]  net821;

wire  [3:0]  slf_op_13_03;

wire  [0:7]  net953;

wire  [0:47]  net826;

wire  [0:47]  net1472;

wire  [3:0]  slf_op_13_05;

wire  [0:47]  net1432;

wire  [0:47]  net1133;

wire  [0:23]  net946;

wire  [0:23]  net825;

wire  [0:47]  net920;

wire  [0:47]  net1226;

wire  [0:23]  net900;

wire  [0:23]  net1378;

wire  [0:47]  net1495;

wire  [0:7]  net1234;

wire  [0:7]  net824;

wire  [0:7]  net861;

wire  [0:47]  net1205;

wire  [0:7]  net1324;

wire  [0:47]  net1292;

wire  [0:7]  net966;

wire  [0:23]  net1335;

wire  [0:23]  net1336;

wire  [0:7]  net860;

wire  [0:23]  net1337;

wire  [0:23]  net1008;

wire  [0:47]  net1158;

wire  [0:23]  net1061;

wire  [0:7]  net1265;

wire  [0:47]  net923;

wire  [0:23]  net829;

wire  [3:0]  slf_op_13_04;

wire  [0:23]  net1059;

wire  [0:23]  net1427;

wire  [0:23]  net1102;

wire  [0:47]  net940;

wire  [0:47]  net1065;

wire  [0:47]  net1015;

wire  [0:47]  net1111;

wire  [0:23]  net1429;

wire  [0:7]  net1325;

wire  [0:23]  net943;

wire  [0:47]  net1249;

wire  [0:7]  net840;

wire  [0:47]  net1157;

wire  [0:47]  net1019;

wire  [0:47]  net1198;

wire  [0:7]  net959;

wire  [0:47]  net1042;

wire  [3:0]  slf_op_10_00;

wire  [3:0]  slf_op_08_00;

wire  [0:7]  net991;

wire  [3:0]  slf_op_13_06;

wire  [0:7]  net999;

wire  [0:47]  net1296;

wire  [0:47]  net822;

wire  [0:47]  net1021;

wire  [0:47]  net1485;

wire  [0:47]  net1020;

wire  [0:23]  net1153;

wire  [0:7]  net1183;

wire  [0:23]  net1010;

wire  [3:0]  slf_op_11_00;

wire  [0:23]  net1011;

wire  [0:23]  net1103;

wire  [0:47]  net1316;

wire  [0:47]  net1066;

wire  [0:47]  net916;

wire  [0:23]  net841;

wire  [0:0]  padinlat_b_r;

wire  [0:7]  net956;

wire  [0:47]  net830;

wire  [0:7]  net1173;

wire  [0:47]  net838;

wire  [0:47]  net1341;

wire  [0:23]  net902;

wire  [0:47]  net921;

wire  [0:23]  net1101;

wire  [0:47]  net1039;

wire  [0:47]  net1247;

wire  [0:47]  net1106;

wire  [0:7]  net1469;

wire  [0:7]  net01070;

wire  [0:47]  net1315;

wire  [3:0]  slf_op_09_00;

wire  [0:47]  net1203;



ice1f_array_RGT_IO_bot9io I_preio_rgt_b13 ( .padin(padin_r_b[8:0]),
     .pado(pado_r_b[8:0]), .padeb(padeb_r_b[8:0]),
     .spi_ss_in_b(spi_ss_in_r[15:0]), .spioeb(spioeb_r[15:0]),
     .spiout(spiout_r[15:0]), .cf_r(cf_r[191:0]),
     .bnl_op_13_01({slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0], slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0]}), .SP4_h_r_13_01(net1481[0:47]),
     .SP4_h_r_13_02(net1495[0:47]), .SP4_h_r_13_03(net1485[0:47]),
     .SP4_h_r_13_04(net1506[0:47]), .SP4_h_r_13_05(net1480[0:47]),
     .SP4_h_r_13_06(net1496[0:47]), .SP4_h_r_13_07(net1472[0:47]),
     .SP4_h_r_13_08(net1407[0:47]), .SP12_h_r_13_01(net1379[0:23]),
     .SP12_h_r_13_02(net1378[0:23]), .SP12_h_r_13_03(net1377[0:23]),
     .SP12_h_r_13_04(net1376[0:23]), .SP12_h_r_13_05(net1426[0:23]),
     .SP12_h_r_13_06(net1427[0:23]), .SP12_h_r_13_07(net1428[0:23]),
     .SP12_h_r_13_08(net1429[0:23]), .rgt_op_13_02(net1175[0:7]),
     .rgt_op_13_03(net1173[0:7]), .rgt_op_13_04(net1183[0:7]),
     .rgt_op_13_05(net1234[0:7]), .rgt_op_13_06(net1233[0:7]),
     .rgt_op_13_07(net1232[0:7]), .rgt_op_13_08(slf_op_12_08[7:0]),
     .slf_op_13_01(slf_op_13_01[3:0]),
     .slf_op_13_02(slf_op_13_02[3:0]),
     .slf_op_13_03(slf_op_13_03[3:0]),
     .slf_op_13_04(slf_op_13_04[3:0]),
     .slf_op_13_05(slf_op_13_05[3:0]),
     .slf_op_13_06(slf_op_13_06[3:0]),
     .slf_op_13_07(slf_op_13_07[3:0]),
     .slf_op_13_08(slf_op_13_08[3:0]),
     .cdone_in(end_of_startup_rgt_b[8:1]),
     .sp4_v_t_13_08(sp4_v_t_13_08[15:0]), .rgt_op_13_01(net840[0:7]),
     .tnl_op_13_08(top_op_12_08[7:0]), .sp4_v_b_13_01(net811[0:15]),
     .wl(wl_r[143:16]), .pgate(pgate_r[143:16]),
     .reset_b(reset_b_r[143:16]), .vdd_cntl(vdd_cntl_r[143:16]),
     .fabric_out_08(net_fabric_out_13_08), .fabric_out_07(net1458),
     .fabric_out_06(net1459), .fabric_out_05(net1461),
     .fabric_out_04(net786), .fabric_out_03(net787),
     .fabric_out_02(net_fabric_out_13_02),
     .fabric_out_01(net_fabric_out_13_01), .shift(shift_br_1),
     .bs_en(bs_en_br_1), .mode(mode_br_1), .sdi(sdio_br_1),
     .hiz_b(hiz_br_1), .prog(prog), .hold(hold_r_b),
     .update(update_br_1), .glb_netwk_col(clk_tree_drv[7:0]),
     .r(r_br_1), .sdo(net800), .bl(bl[329:312]), .tclk(tck_br_1),
     .ceb(ceb_br_1));
ice1f_array_BOT_IO_rgt12io I_preio_bot_r ( .padin_b_r(padin_b_r[11:0]),
     .padeb_b_r(padeb_b_r[11:0]), .pado_b_r(pado_b_r[11:0]),
     .spiceb(spioeb[11:0]), .spiout(spiout[11:0]),
     .spi_ss_in_b(spi_ss_in_b[11:0]), .tnr_op_06_00({slf_op_13_01[3],
     slf_op_13_01[2], slf_op_13_01[1], slf_op_13_01[0],
     slf_op_13_01[3], slf_op_13_01[2], slf_op_13_01[1],
     slf_op_13_01[0]}), .sp4_h_r_06_00(net811[0:15]),
     .fabric_out_12_00(net_fabric_out_12_00),
     .end_of_startup_top_l(end_of_startup_bot_r[12:7]),
     .cf_bot_r(cf_b[143:0]), .fabric_out_07_00(net_fabric_out_07_00),
     .bl_04(bl[203:162]), .bnl_op_01_00(rgt_op_07_01[7:0]),
     .sp4_v_b_01_00(sp4_v_b_07_01[47:0]),
     .slf_op_01_00(slf_op_07_00[3:0]),
     .lft_op_01_00(slf_op_07_01[7:0]), .sp12_v_b_01_00(net821[0:23]),
     .sp4_v_b_02_00(net822[0:47]), .slf_op_02_00(slf_op_08_00[3:0]),
     .lft_op_02_00(net824[0:7]), .sp12_v_b_02_00(net825[0:23]),
     .sp4_v_b_03_00(net826[0:47]), .slf_op_03_00(slf_op_09_00[3:0]),
     .lft_op_03_00(net828[0:7]), .sp12_v_b_03_00(net829[0:23]),
     .sp4_v_b_04_00(net830[0:47]), .slf_op_04_00(slf_op_10_00[3:0]),
     .lft_op_04_00(net1493[0:7]), .sp12_v_b_04_00(net833[0:23]),
     .sp4_v_b_05_00(net834[0:47]), .slf_op_05_00(slf_op_11_00[3:0]),
     .lft_op_05_00(net836[0:7]), .sp12_v_b_05_00(net837[0:23]),
     .sp4_v_b_06_00(net838[0:47]), .slf_op_06_00(slf_op_12_00[3:0]),
     .lft_op_06_00(net840[0:7]), .sp12_v_b_06_00(net841[0:23]),
     .sp4_h_l_21_00(sp4_h_l_07_00[15:0]), .hold_b_r(hold_b_r),
     .wl_l({wl_r[1], wl_r[0], wl_r[2], wl_r[3], wl_r[5], wl_r[4],
     wl_r[6], wl_r[7], wl_r[9], wl_r[8], wl_r[10], wl_r[11], wl_r[13],
     wl_r[12], wl_r[14], wl_r[15]}), .vdd_cntl_l({vdd_cntl_r[1],
     vdd_cntl_r[0], vdd_cntl_r[2], vdd_cntl_r[3], vdd_cntl_r[5],
     vdd_cntl_r[4], vdd_cntl_r[6], vdd_cntl_r[7], vdd_cntl_r[9],
     vdd_cntl_r[8], vdd_cntl_r[10], vdd_cntl_r[11], vdd_cntl_r[13],
     vdd_cntl_r[12], vdd_cntl_r[14], vdd_cntl_r[15]}),
     .update_i(update_i), .tclk_i(tclk_i), .shift_i(shift_i),
     .sdi(sdi), .reset_l({reset_b_r[1], reset_b_r[0], reset_b_r[2],
     reset_b_r[3], reset_b_r[5], reset_b_r[4], reset_b_r[6],
     reset_b_r[7], reset_b_r[9], reset_b_r[8], reset_b_r[10],
     reset_b_r[11], reset_b_r[13], reset_b_r[12], reset_b_r[14],
     reset_b_r[15]}), .r_i(r_i), .prog(prog), .pgate_l({pgate_r[1],
     pgate_r[0], pgate_r[2], pgate_r[3], pgate_r[5], pgate_r[4],
     pgate_r[6], pgate_r[7], pgate_r[9], pgate_r[8], pgate_r[10],
     pgate_r[11], pgate_r[13], pgate_r[12], pgate_r[14], pgate_r[15]}),
     .mode_i(mode_i), .hiz_b_i(hiz_b_i), .bs_en_i(bs_en_i),
     .sdo(sdo_pad), .glb_net_06(net0855[0:7]),
     .glb_net_05(net0856[0:7]), .glb_net_04(net860[0:7]),
     .glb_net_03(net861[0:7]), .glb_net_02(net0859[0:7]),
     .glb_net_01(net0860[0:7]), .bl_06(bl[311:258]),
     .bl_05(bl[257:204]), .bl_03(bl[161:108]), .bl_02(bl[107:54]),
     .bl_01(bl[53:0]), .ceb_i(ceb_i));
pinlatbuf12p I_pinlatbuf12p_b ( .pad_in(padin_b_r[0]),
     .icegate(hold_b_r), .cbit(cf_b[15]), .cout(padinlat_b_r[0]),
     .prog(prog));
pinlatbuf12p I_pinlatbuf12p ( .pad_in(padin_r_b[8]),
     .icegate(hold_r_b), .cbit(cf_r[183]), .cout(padinlat_r_b[11]),
     .prog(prog));
scanbuf1f I_scanbuf_mr ( .update_i(update_br_1), .tclk_i(tck_br_1),
     .shift_i(shift_br_1), .sdi(net800), .r_i(r_br_1),
     .mode_i(mode_br_1), .hiz_b_i(hiz_br_1), .ceb_i(ceb_br_1),
     .bs_en_i(bs_en_br_1), .update_o(update_o), .tclk_o(tclk_o),
     .shift_o(shift_o), .sdo(sdo), .r_o(r_o), .mode_o(mode_o),
     .hiz_b_o(hiz_b_o), .ceb_o(ceb_o), .bs_en_o(bs_en_o));
scanbuf1f I_scanbuf_br0 ( .update_i(update_mi), .tclk_i(tclk_mi),
     .shift_i(shift_mi), .sdi(sdi_pad), .r_i(r_mi), .mode_i(mode_mi),
     .hiz_b_i(hiz_b_mi), .ceb_i(ceb_mi), .bs_en_i(bs_en_mi),
     .update_o(update_br_1), .tclk_o(tck_br_1), .shift_o(shift_br_1),
     .sdo(sdio_br_1), .r_o(r_br_1), .mode_o(mode_br_1),
     .hiz_b_o(hiz_br_1), .ceb_o(ceb_br_1), .bs_en_o(bs_en_br_1));
ice1f_array_BRAM_bot I_bram_col_b10 ( .glb_netwk_top(net1469[0:7]),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .vdd_cntl(vdd_cntl_r[143:16]), .wl(wl_r[143:16]),
     .sp12_v_t_08(sp12_v_t_10_08[23:0]), .top_op_08(top_op_10_08[7:0]),
     .sp4_v_t_08(sp4_v_t_10_08[47:0]), .tnl_op_08(tnl_op_10_08[7:0]),
     .tnr_op_08(tnr_op_10_08[7:0]), .glb_netwk_bot(net860[0:7]),
     .bm_init_i(bm_init_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sweb_i(bm_sweb_i[1:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sdi_i(bm_sdi_i[1:0]),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sweb_o(bm_sweb_o[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .prog(prog),
     .glb_netwk_col(clk_tree_drv[7:0]), .sp12_h_l_07(net1152[0:23]),
     .sp4_v_b_08(net1158[0:47]), .bnr_op_01({slf_op_11_00[3],
     slf_op_11_00[2], slf_op_11_00[1], slf_op_11_00[0],
     slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0]}), .sp12_h_r_06(net900[0:23]),
     .sp12_h_l_06(net1151[0:23]), .sp12_h_r_05(net902[0:23]),
     .sp12_h_r_08(net903[0:23]), .sp12_h_r_03(net904[0:23]),
     .sp12_h_l_08(net1153[0:23]), .sp12_h_l_05(net1150[0:23]),
     .sp12_h_r_07(net907[0:23]), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_sreb_o(bm_sreb_o), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .sp4_r_v_b_01(net834[0:47]),
     .sp4_v_b_02(net1108[0:47]), .sp4_r_v_b_02(net916[0:47]),
     .sp4_v_b_03(net1107[0:47]), .sp4_r_v_b_03(net918[0:47]),
     .sp4_v_b_04(net1106[0:47]), .sp4_r_v_b_04(net920[0:47]),
     .sp4_r_v_b_06(net921[0:47]), .sp4_v_b_06(net1156[0:47]),
     .sp4_r_v_b_05(net923[0:47]), .sp4_v_b_05(net1155[0:47]),
     .lft_op_08(slf_op_09_08[7:0]), .lft_op_07(net1324[0:7]),
     .lft_op_06(net1325[0:7]), .lft_op_05(net1326[0:7]),
     .sp4_v_b_07(net1157[0:47]), .sp12_h_l_03(net1101[0:23]),
     .sp12_h_l_04(net1100[0:23]), .sp12_h_l_02(net1102[0:23]),
     .sp12_h_l_01(net1103[0:23]), .slf_op_07(net1140[0:7]),
     .slf_op_08(slf_op_10_08[7:0]), .sp4_h_l_07(net1132[0:47]),
     .sp4_h_l_08(net1131[0:47]), .sp4_h_r_07(net938[0:47]),
     .sp4_h_r_08(net939[0:47]), .sp4_r_v_b_07(net940[0:47]),
     .sp4_r_v_b_08(net941[0:47]), .sp4_v_b_01(net830[0:47]),
     .sp12_h_r_01(net943[0:23]), .sp12_h_r_02(net944[0:23]),
     .bl(bl[203:162]), .sp12_h_r_04(net946[0:23]),
     .sp12_v_b_01(net833[0:23]), .bnl_op_01({slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0],
     slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0]}), .lft_op_01(net828[0:7]),
     .lft_op_02(net1267[0:7]), .lft_op_03(net1265[0:7]),
     .lft_op_04(net1275[0:7]), .rgt_op_07(net953[0:7]),
     .rgt_op_08(slf_op_11_08[7:0]), .bot_op_01({slf_op_10_00[3],
     slf_op_10_00[2], slf_op_10_00[1], slf_op_10_00[0],
     slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0]}), .rgt_op_03(net956[0:7]),
     .rgt_op_02(net957[0:7]), .rgt_op_01(net836[0:7]),
     .rgt_op_04(net959[0:7]), .slf_op_04(net1091[0:7]),
     .slf_op_03(net1081[0:7]), .slf_op_02(net1083[0:7]),
     .slf_op_01(net1493[0:7]), .slf_op_06(net1141[0:7]),
     .rgt_op_05(net965[0:7]), .rgt_op_06(net966[0:7]),
     .slf_op_05(net1142[0:7]), .sp4_h_r_04(net968[0:47]),
     .sp4_h_r_03(net969[0:47]), .sp4_h_r_02(net970[0:47]),
     .sp4_h_r_01(net971[0:47]), .sp4_h_l_04(net1110[0:47]),
     .sp4_h_l_03(net1111[0:47]), .sp4_h_l_02(net1112[0:47]),
     .sp4_h_l_01(net1113[0:47]), .sp4_h_r_06(net976[0:47]),
     .sp4_h_l_06(net1133[0:47]), .sp4_h_r_05(net978[0:47]),
     .sp4_h_l_05(net1134[0:47]));
ice1f_array_LT_top I_lt_col_b07 ( .glb_netwk_to(net863[0:7]),
     .glb_netwk_bo(net0860[0:7]), .vdd_cntl(vdd_cntl_r[143:16]),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .top_op_08(top_op_07_08[7:0]), .tnl_op_08(tnl_op_07_08[7:0]),
     .tnr_op_08(tnr_op_07_08[7:0]), .sp12_v_t_08(sp12_v_t_07_08[23:0]),
     .sp4_v_t_08(sp4_v_t_07_08[47:0]), .wl(wl_r[143:16]),
     .rgt_op_03(net989[0:7]), .slf_op_02(slf_op_07_02[7:0]),
     .rgt_op_02(net991[0:7]), .rgt_op_01(net824[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(rgt_op_07_04[7:0]),
     .lft_op_03(rgt_op_07_03[7:0]), .lft_op_02(rgt_op_07_02[7:0]),
     .lft_op_01(rgt_op_07_01[7:0]), .rgt_op_04(net999[0:7]),
     .carry_in(net1462), .bnl_op_01({bnl_op_07_01[3], bnl_op_07_01[2],
     bnl_op_07_01[1], bnl_op_07_01[0], bnl_op_07_01[3],
     bnl_op_07_01[2], bnl_op_07_01[1], bnl_op_07_01[0]}),
     .slf_op_04(slf_op_07_04[7:0]), .slf_op_03(slf_op_07_03[7:0]),
     .slf_op_01(slf_op_07_01[7:0]), .sp4_h_l_04(sp4_h_l_07_04[47:0]),
     .carry_out(carry_out_07_08), .sp12_v_b__01(net821[0:23]),
     .sp12_h_r_04(net1008[0:23]), .sp12_h_r_03(net1009[0:23]),
     .sp12_h_r_02(net1010[0:23]), .sp12_h_r_01(net1011[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_07_01[47:0]), .sp4_r_v_b_04(net1014[0:47]),
     .sp4_r_v_b_03(net1015[0:47]), .sp4_r_v_b_02(net1016[0:47]),
     .sp4_r_v_b_01(net822[0:47]), .sp4_h_r_04(net1018[0:47]),
     .sp4_h_r_03(net1019[0:47]), .sp4_h_r_02(net1020[0:47]),
     .sp4_h_r_01(net1021[0:47]), .sp4_h_l_03(sp4_h_l_07_03[47:0]),
     .sp4_h_l_02(sp4_h_l_07_02[47:0]),
     .sp4_h_l_01(sp4_h_l_07_01[47:0]), .bl(bl[53:0]),
     .bot_op_01({slf_op_07_00[3], slf_op_07_00[2], slf_op_07_00[1],
     slf_op_07_00[0], slf_op_07_00[3], slf_op_07_00[2],
     slf_op_07_00[1], slf_op_07_00[0]}),
     .sp12_h_l_01(sp12_h_l_07_01[23:0]),
     .sp12_h_l_02(sp12_h_l_07_02[23:0]),
     .sp12_h_l_03(sp12_h_l_07_03[23:0]),
     .sp12_h_l_04(sp12_h_l_07_04[23:0]),
     .sp4_v_b_04(sp4_v_b_07_04[47:0]),
     .sp4_v_b_03(sp4_v_b_07_03[47:0]),
     .sp4_v_b_02(sp4_v_b_07_02[47:0]), .bnr_op_01({slf_op_08_00[3],
     slf_op_08_00[2], slf_op_08_00[1], slf_op_08_00[0],
     slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0]}), .sp4_h_l_05(sp4_h_l_07_05[47:0]),
     .sp4_h_l_06(sp4_h_l_07_06[47:0]),
     .sp4_h_l_07(sp4_h_l_07_07[47:0]),
     .sp4_h_l_08(sp4_h_l_07_08[47:0]), .sp4_h_r_08(net1039[0:47]),
     .sp4_h_r_07(net1040[0:47]), .sp4_h_r_06(net1041[0:47]),
     .sp4_h_r_05(net1042[0:47]), .slf_op_05(slf_op_07_05[7:0]),
     .slf_op_06(slf_op_07_06[7:0]), .slf_op_07(slf_op_07_07[7:0]),
     .slf_op_08(slf_op_07_08[7:0]), .rgt_op_08(slf_op_08_08[7:0]),
     .rgt_op_07(net1048[0:7]), .rgt_op_06(net1049[0:7]),
     .rgt_op_05(net1050[0:7]), .lft_op_08(rgt_op_07_08[7:0]),
     .lft_op_07(rgt_op_07_07[7:0]), .lft_op_06(rgt_op_07_06[7:0]),
     .lft_op_05(rgt_op_07_05[7:0]), .sp12_h_l_08(sp12_h_l_07_08[23:0]),
     .sp12_h_l_07(sp12_h_l_07_07[23:0]),
     .sp12_h_l_06(sp12_h_l_07_06[23:0]), .sp12_h_r_05(net1058[0:23]),
     .sp12_h_r_06(net1059[0:23]), .sp12_h_r_07(net1060[0:23]),
     .sp12_h_r_08(net1061[0:23]), .sp12_h_l_05(sp12_h_l_07_05[23:0]),
     .sp4_r_v_b_05(net1063[0:47]), .sp4_r_v_b_06(net1064[0:47]),
     .sp4_r_v_b_07(net1065[0:47]), .sp4_r_v_b_08(net1066[0:47]),
     .sp4_v_b_08(sp4_v_b_07_08[47:0]),
     .sp4_v_b_07(sp4_v_b_07_07[47:0]),
     .sp4_v_b_06(sp4_v_b_07_06[47:0]),
     .sp4_v_b_05(sp4_v_b_07_05[47:0]));
ice1f_array_LT_top I_lt_col_b09 ( .glb_netwk_to(net01070[0:7]),
     .glb_netwk_bo(net861[0:7]), .vdd_cntl(vdd_cntl_r[143:16]),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .top_op_08(top_op_09_08[7:0]), .tnl_op_08(tnl_op_09_08[7:0]),
     .tnr_op_08(tnr_op_09_08[7:0]), .sp12_v_t_08(sp12_v_t_09_08[23:0]),
     .sp4_v_t_08(sp4_v_t_09_08[47:0]), .wl(wl_r[143:16]),
     .rgt_op_03(net1081[0:7]), .slf_op_02(net1267[0:7]),
     .rgt_op_02(net1083[0:7]), .rgt_op_01(net1493[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net999[0:7]), .lft_op_03(net989[0:7]),
     .lft_op_02(net991[0:7]), .lft_op_01(net824[0:7]),
     .rgt_op_04(net1091[0:7]), .carry_in(net1092),
     .bnl_op_01({slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0], slf_op_08_00[3], slf_op_08_00[2],
     slf_op_08_00[1], slf_op_08_00[0]}), .slf_op_04(net1275[0:7]),
     .slf_op_03(net1265[0:7]), .slf_op_01(net828[0:7]),
     .sp4_h_l_04(net1294[0:47]), .carry_out(carry_out_09_08),
     .sp12_v_b__01(net829[0:23]), .sp12_h_r_04(net1100[0:23]),
     .sp12_h_r_03(net1101[0:23]), .sp12_h_r_02(net1102[0:23]),
     .sp12_h_r_01(net1103[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(net826[0:47]), .sp4_r_v_b_04(net1106[0:47]),
     .sp4_r_v_b_03(net1107[0:47]), .sp4_r_v_b_02(net1108[0:47]),
     .sp4_r_v_b_01(net830[0:47]), .sp4_h_r_04(net1110[0:47]),
     .sp4_h_r_03(net1111[0:47]), .sp4_h_r_02(net1112[0:47]),
     .sp4_h_r_01(net1113[0:47]), .sp4_h_l_03(net1295[0:47]),
     .sp4_h_l_02(net1296[0:47]), .sp4_h_l_01(net1297[0:47]),
     .bl(bl[161:108]), .bot_op_01({slf_op_09_00[3], slf_op_09_00[2],
     slf_op_09_00[1], slf_op_09_00[0], slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0]}),
     .sp12_h_l_01(net1287[0:23]), .sp12_h_l_02(net1286[0:23]),
     .sp12_h_l_03(net1285[0:23]), .sp12_h_l_04(net1284[0:23]),
     .sp4_v_b_04(net1290[0:47]), .sp4_v_b_03(net1291[0:47]),
     .sp4_v_b_02(net1292[0:47]), .bnr_op_01({slf_op_10_00[3],
     slf_op_10_00[2], slf_op_10_00[1], slf_op_10_00[0],
     slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0]}), .sp4_h_l_05(net1318[0:47]),
     .sp4_h_l_06(net1317[0:47]), .sp4_h_l_07(net1316[0:47]),
     .sp4_h_l_08(net1315[0:47]), .sp4_h_r_08(net1131[0:47]),
     .sp4_h_r_07(net1132[0:47]), .sp4_h_r_06(net1133[0:47]),
     .sp4_h_r_05(net1134[0:47]), .slf_op_05(net1326[0:7]),
     .slf_op_06(net1325[0:7]), .slf_op_07(net1324[0:7]),
     .slf_op_08(slf_op_09_08[7:0]), .rgt_op_08(slf_op_10_08[7:0]),
     .rgt_op_07(net1140[0:7]), .rgt_op_06(net1141[0:7]),
     .rgt_op_05(net1142[0:7]), .lft_op_08(slf_op_08_08[7:0]),
     .lft_op_07(net1048[0:7]), .lft_op_06(net1049[0:7]),
     .lft_op_05(net1050[0:7]), .sp12_h_l_08(net1337[0:23]),
     .sp12_h_l_07(net1336[0:23]), .sp12_h_l_06(net1335[0:23]),
     .sp12_h_r_05(net1150[0:23]), .sp12_h_r_06(net1151[0:23]),
     .sp12_h_r_07(net1152[0:23]), .sp12_h_r_08(net1153[0:23]),
     .sp12_h_l_05(net1334[0:23]), .sp4_r_v_b_05(net1155[0:47]),
     .sp4_r_v_b_06(net1156[0:47]), .sp4_r_v_b_07(net1157[0:47]),
     .sp4_r_v_b_08(net1158[0:47]), .sp4_v_b_08(net1342[0:47]),
     .sp4_v_b_07(net1341[0:47]), .sp4_v_b_06(net1340[0:47]),
     .sp4_v_b_05(net1339[0:47]));
ice1f_array_LT_top I_lt_col_b11 ( .glb_netwk_to(net859[0:7]),
     .glb_netwk_bo(net0856[0:7]), .vdd_cntl(vdd_cntl_r[143:16]),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .top_op_08(top_op_11_08[7:0]), .tnl_op_08(tnl_op_11_08[7:0]),
     .tnr_op_08(tnr_op_11_08[7:0]), .sp12_v_t_08(sp12_v_t_11_08[23:0]),
     .sp4_v_t_08(sp4_v_t_11_08[47:0]), .wl(wl_r[143:16]),
     .rgt_op_03(net1173[0:7]), .slf_op_02(net957[0:7]),
     .rgt_op_02(net1175[0:7]), .rgt_op_01(net840[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net1091[0:7]), .lft_op_03(net1081[0:7]),
     .lft_op_02(net1083[0:7]), .lft_op_01(net1493[0:7]),
     .rgt_op_04(net1183[0:7]), .carry_in(net1507),
     .bnl_op_01({slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0], slf_op_10_00[3], slf_op_10_00[2],
     slf_op_10_00[1], slf_op_10_00[0]}), .slf_op_04(net959[0:7]),
     .slf_op_03(net956[0:7]), .slf_op_01(net836[0:7]),
     .sp4_h_l_04(net968[0:47]), .carry_out(carry_out_11_08),
     .sp12_v_b__01(net837[0:23]), .sp12_h_r_04(net1192[0:23]),
     .sp12_h_r_03(net1193[0:23]), .sp12_h_r_02(net1194[0:23]),
     .sp12_h_r_01(net1195[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(net834[0:47]), .sp4_r_v_b_04(net1198[0:47]),
     .sp4_r_v_b_03(net1199[0:47]), .sp4_r_v_b_02(net1200[0:47]),
     .sp4_r_v_b_01(net838[0:47]), .sp4_h_r_04(net1202[0:47]),
     .sp4_h_r_03(net1203[0:47]), .sp4_h_r_02(net1204[0:47]),
     .sp4_h_r_01(net1205[0:47]), .sp4_h_l_03(net969[0:47]),
     .sp4_h_l_02(net970[0:47]), .sp4_h_l_01(net971[0:47]),
     .bl(bl[257:204]), .bot_op_01({slf_op_11_00[3], slf_op_11_00[2],
     slf_op_11_00[1], slf_op_11_00[0], slf_op_11_00[3],
     slf_op_11_00[2], slf_op_11_00[1], slf_op_11_00[0]}),
     .sp12_h_l_01(net943[0:23]), .sp12_h_l_02(net944[0:23]),
     .sp12_h_l_03(net904[0:23]), .sp12_h_l_04(net946[0:23]),
     .sp4_v_b_04(net920[0:47]), .sp4_v_b_03(net918[0:47]),
     .sp4_v_b_02(net916[0:47]), .bnr_op_01({slf_op_12_00[3],
     slf_op_12_00[2], slf_op_12_00[1], slf_op_12_00[0],
     slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0]}), .sp4_h_l_05(net978[0:47]),
     .sp4_h_l_06(net976[0:47]), .sp4_h_l_07(net938[0:47]),
     .sp4_h_l_08(net939[0:47]), .sp4_h_r_08(net1223[0:47]),
     .sp4_h_r_07(net1224[0:47]), .sp4_h_r_06(net1225[0:47]),
     .sp4_h_r_05(net1226[0:47]), .slf_op_05(net965[0:7]),
     .slf_op_06(net966[0:7]), .slf_op_07(net953[0:7]),
     .slf_op_08(slf_op_11_08[7:0]), .rgt_op_08(slf_op_12_08[7:0]),
     .rgt_op_07(net1232[0:7]), .rgt_op_06(net1233[0:7]),
     .rgt_op_05(net1234[0:7]), .lft_op_08(slf_op_10_08[7:0]),
     .lft_op_07(net1140[0:7]), .lft_op_06(net1141[0:7]),
     .lft_op_05(net1142[0:7]), .sp12_h_l_08(net903[0:23]),
     .sp12_h_l_07(net907[0:23]), .sp12_h_l_06(net900[0:23]),
     .sp12_h_r_05(net1242[0:23]), .sp12_h_r_06(net1243[0:23]),
     .sp12_h_r_07(net1244[0:23]), .sp12_h_r_08(net1245[0:23]),
     .sp12_h_l_05(net902[0:23]), .sp4_r_v_b_05(net1247[0:47]),
     .sp4_r_v_b_06(net1248[0:47]), .sp4_r_v_b_07(net1249[0:47]),
     .sp4_r_v_b_08(net1250[0:47]), .sp4_v_b_08(net941[0:47]),
     .sp4_v_b_07(net940[0:47]), .sp4_v_b_06(net921[0:47]),
     .sp4_v_b_05(net923[0:47]));
ice1f_array_LT_top I_lt_col_b08 ( .glb_netwk_to(net862[0:7]),
     .glb_netwk_bo(net0859[0:7]), .vdd_cntl(vdd_cntl_r[143:16]),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .top_op_08(top_op_08_08[7:0]), .tnl_op_08(tnl_op_08_08[7:0]),
     .tnr_op_08(tnr_op_08_08[7:0]), .sp12_v_t_08(sp12_v_t_08_08[23:0]),
     .sp4_v_t_08(sp4_v_t_08_08[47:0]), .wl(wl_r[143:16]),
     .rgt_op_03(net1265[0:7]), .slf_op_02(net991[0:7]),
     .rgt_op_02(net1267[0:7]), .rgt_op_01(net828[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(slf_op_07_04[7:0]),
     .lft_op_03(slf_op_07_03[7:0]), .lft_op_02(slf_op_07_02[7:0]),
     .lft_op_01(slf_op_07_01[7:0]), .rgt_op_04(net1275[0:7]),
     .carry_in(net1276), .bnl_op_01({slf_op_07_00[3], slf_op_07_00[2],
     slf_op_07_00[1], slf_op_07_00[0], slf_op_07_00[3],
     slf_op_07_00[2], slf_op_07_00[1], slf_op_07_00[0]}),
     .slf_op_04(net999[0:7]), .slf_op_03(net989[0:7]),
     .slf_op_01(net824[0:7]), .sp4_h_l_04(net1018[0:47]),
     .carry_out(carry_out_08_08), .sp12_v_b__01(net825[0:23]),
     .sp12_h_r_04(net1284[0:23]), .sp12_h_r_03(net1285[0:23]),
     .sp12_h_r_02(net1286[0:23]), .sp12_h_r_01(net1287[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .sp4_v_b_01(net822[0:47]),
     .sp4_r_v_b_04(net1290[0:47]), .sp4_r_v_b_03(net1291[0:47]),
     .sp4_r_v_b_02(net1292[0:47]), .sp4_r_v_b_01(net826[0:47]),
     .sp4_h_r_04(net1294[0:47]), .sp4_h_r_03(net1295[0:47]),
     .sp4_h_r_02(net1296[0:47]), .sp4_h_r_01(net1297[0:47]),
     .sp4_h_l_03(net1019[0:47]), .sp4_h_l_02(net1020[0:47]),
     .sp4_h_l_01(net1021[0:47]), .bl(bl[107:54]),
     .bot_op_01({slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0], slf_op_08_00[3], slf_op_08_00[2],
     slf_op_08_00[1], slf_op_08_00[0]}), .sp12_h_l_01(net1011[0:23]),
     .sp12_h_l_02(net1010[0:23]), .sp12_h_l_03(net1009[0:23]),
     .sp12_h_l_04(net1008[0:23]), .sp4_v_b_04(net1014[0:47]),
     .sp4_v_b_03(net1015[0:47]), .sp4_v_b_02(net1016[0:47]),
     .bnr_op_01({slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0], slf_op_09_00[3], slf_op_09_00[2],
     slf_op_09_00[1], slf_op_09_00[0]}), .sp4_h_l_05(net1042[0:47]),
     .sp4_h_l_06(net1041[0:47]), .sp4_h_l_07(net1040[0:47]),
     .sp4_h_l_08(net1039[0:47]), .sp4_h_r_08(net1315[0:47]),
     .sp4_h_r_07(net1316[0:47]), .sp4_h_r_06(net1317[0:47]),
     .sp4_h_r_05(net1318[0:47]), .slf_op_05(net1050[0:7]),
     .slf_op_06(net1049[0:7]), .slf_op_07(net1048[0:7]),
     .slf_op_08(slf_op_08_08[7:0]), .rgt_op_08(slf_op_09_08[7:0]),
     .rgt_op_07(net1324[0:7]), .rgt_op_06(net1325[0:7]),
     .rgt_op_05(net1326[0:7]), .lft_op_08(slf_op_07_08[7:0]),
     .lft_op_07(slf_op_07_07[7:0]), .lft_op_06(slf_op_07_06[7:0]),
     .lft_op_05(slf_op_07_05[7:0]), .sp12_h_l_08(net1061[0:23]),
     .sp12_h_l_07(net1060[0:23]), .sp12_h_l_06(net1059[0:23]),
     .sp12_h_r_05(net1334[0:23]), .sp12_h_r_06(net1335[0:23]),
     .sp12_h_r_07(net1336[0:23]), .sp12_h_r_08(net1337[0:23]),
     .sp12_h_l_05(net1058[0:23]), .sp4_r_v_b_05(net1339[0:47]),
     .sp4_r_v_b_06(net1340[0:47]), .sp4_r_v_b_07(net1341[0:47]),
     .sp4_r_v_b_08(net1342[0:47]), .sp4_v_b_08(net1066[0:47]),
     .sp4_v_b_07(net1065[0:47]), .sp4_v_b_06(net1064[0:47]),
     .sp4_v_b_05(net1063[0:47]));
ice1f_array_LT_top I_lt_col_b12 ( .glb_netwk_to(net858[0:7]),
     .glb_netwk_bo(net0855[0:7]), .vdd_cntl(vdd_cntl_r[143:16]),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .top_op_08(top_op_12_08[7:0]), .tnl_op_08(tnl_op_12_08[7:0]),
     .tnr_op_08(tnr_op_12_08[7:0]), .sp12_v_t_08(sp12_v_t_12_08[23:0]),
     .sp4_v_t_08(sp4_v_t_12_08[47:0]), .wl(wl_r[143:16]),
     .rgt_op_03({slf_op_13_03[3], slf_op_13_03[2], slf_op_13_03[1],
     slf_op_13_03[0], slf_op_13_03[3], slf_op_13_03[2],
     slf_op_13_03[1], slf_op_13_03[0]}), .slf_op_02(net1175[0:7]),
     .rgt_op_02({slf_op_13_02[3], slf_op_13_02[2], slf_op_13_02[1],
     slf_op_13_02[0], slf_op_13_02[3], slf_op_13_02[2],
     slf_op_13_02[1], slf_op_13_02[0]}), .rgt_op_01({slf_op_13_01[3],
     slf_op_13_01[2], slf_op_13_01[1], slf_op_13_01[0],
     slf_op_13_01[3], slf_op_13_01[2], slf_op_13_01[1],
     slf_op_13_01[0]}), .purst(purst), .prog(prog),
     .lft_op_04(net959[0:7]), .lft_op_03(net956[0:7]),
     .lft_op_02(net957[0:7]), .lft_op_01(net836[0:7]),
     .rgt_op_04({slf_op_13_04[3], slf_op_13_04[2], slf_op_13_04[1],
     slf_op_13_04[0], slf_op_13_04[3], slf_op_13_04[2],
     slf_op_13_04[1], slf_op_13_04[0]}), .carry_in(net1368),
     .bnl_op_01({slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0], slf_op_11_00[3], slf_op_11_00[2],
     slf_op_11_00[1], slf_op_11_00[0]}), .slf_op_04(net1183[0:7]),
     .slf_op_03(net1173[0:7]), .slf_op_01(net840[0:7]),
     .sp4_h_l_04(net1202[0:47]), .carry_out(carry_out_12_08),
     .sp12_v_b__01(net841[0:23]), .sp12_h_r_04(net1376[0:23]),
     .sp12_h_r_03(net1377[0:23]), .sp12_h_r_02(net1378[0:23]),
     .sp12_h_r_01(net1379[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(net838[0:47]), .sp4_r_v_b_04(net1382[0:47]),
     .sp4_r_v_b_03(net1383[0:47]), .sp4_r_v_b_02(net1384[0:47]),
     .sp4_r_v_b_01(net1385[0:47]), .sp4_h_r_04(net1506[0:47]),
     .sp4_h_r_03(net1485[0:47]), .sp4_h_r_02(net1495[0:47]),
     .sp4_h_r_01(net1481[0:47]), .sp4_h_l_03(net1203[0:47]),
     .sp4_h_l_02(net1204[0:47]), .sp4_h_l_01(net1205[0:47]),
     .bl(bl[311:258]), .bot_op_01({slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0], slf_op_12_00[3],
     slf_op_12_00[2], slf_op_12_00[1], slf_op_12_00[0]}),
     .sp12_h_l_01(net1195[0:23]), .sp12_h_l_02(net1194[0:23]),
     .sp12_h_l_03(net1193[0:23]), .sp12_h_l_04(net1192[0:23]),
     .sp4_v_b_04(net1198[0:47]), .sp4_v_b_03(net1199[0:47]),
     .sp4_v_b_02(net1200[0:47]), .bnr_op_01({tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .sp4_h_l_05(net1226[0:47]), .sp4_h_l_06(net1225[0:47]),
     .sp4_h_l_07(net1224[0:47]), .sp4_h_l_08(net1223[0:47]),
     .sp4_h_r_08(net1407[0:47]), .sp4_h_r_07(net1472[0:47]),
     .sp4_h_r_06(net1496[0:47]), .sp4_h_r_05(net1480[0:47]),
     .slf_op_05(net1234[0:7]), .slf_op_06(net1233[0:7]),
     .slf_op_07(net1232[0:7]), .slf_op_08(slf_op_12_08[7:0]),
     .rgt_op_08({slf_op_13_08[3], slf_op_13_08[2], slf_op_13_08[1],
     slf_op_13_08[0], slf_op_13_08[3], slf_op_13_08[2],
     slf_op_13_08[1], slf_op_13_08[0]}), .rgt_op_07({slf_op_13_07[3],
     slf_op_13_07[2], slf_op_13_07[1], slf_op_13_07[0],
     slf_op_13_07[3], slf_op_13_07[2], slf_op_13_07[1],
     slf_op_13_07[0]}), .rgt_op_06({slf_op_13_06[3], slf_op_13_06[2],
     slf_op_13_06[1], slf_op_13_06[0], slf_op_13_06[3],
     slf_op_13_06[2], slf_op_13_06[1], slf_op_13_06[0]}),
     .rgt_op_05({slf_op_13_05[3], slf_op_13_05[2], slf_op_13_05[1],
     slf_op_13_05[0], slf_op_13_05[3], slf_op_13_05[2],
     slf_op_13_05[1], slf_op_13_05[0]}), .lft_op_08(slf_op_11_08[7:0]),
     .lft_op_07(net953[0:7]), .lft_op_06(net966[0:7]),
     .lft_op_05(net965[0:7]), .sp12_h_l_08(net1245[0:23]),
     .sp12_h_l_07(net1244[0:23]), .sp12_h_l_06(net1243[0:23]),
     .sp12_h_r_05(net1426[0:23]), .sp12_h_r_06(net1427[0:23]),
     .sp12_h_r_07(net1428[0:23]), .sp12_h_r_08(net1429[0:23]),
     .sp12_h_l_05(net1242[0:23]), .sp4_r_v_b_05(net1431[0:47]),
     .sp4_r_v_b_06(net1432[0:47]), .sp4_r_v_b_07(net1433[0:47]),
     .sp4_r_v_b_08(net1434[0:47]), .sp4_v_b_08(net1250[0:47]),
     .sp4_v_b_07(net1249[0:47]), .sp4_v_b_06(net1248[0:47]),
     .sp4_v_b_05(net1247[0:47]));
fabric_outbuf12p I_fbuf_2 ( .fabric_out(net_fabric_out_13_02),
     .cout(fabric_out_13_02));
fabric_outbuf12p I_fbuf_5 ( .fabric_out(padinlat_b_r[0]),
     .cout(padin_07_00a));
fabric_outbuf12p I_fbuf_1 ( .fabric_out(net_fabric_out_13_08),
     .cout(fabric_out_13_08));
fabric_outbuf12p I_fbuf_0 ( .fabric_out(padinlat_r_b[11]),
     .cout(padin_13_08b));
fabric_outbuf12p I_fbuf_4 ( .fabric_out(net_fabric_out_12_00),
     .cout(fabric_out_12_00));
fabric_outbuf12p I_fbuf_3 ( .fabric_out(net_fabric_out_13_01),
     .cout(fabric_out_13_01));
fabric_outbuf12p I_fbuf_7 ( .fabric_out(net_fabric_out_07_00),
     .cout(fabric_out_07_00));
clk_quad_buf12px8 I_clk_quadbuf12px8 ( .clko(clk_tree_drv[7:0]),
     .clki(glb_in[7:0]));

endmodule
// Library - misc, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:59 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_mux2_hvt ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - leafcell, Cell - ice1f_array_RGT_IO_top12io, View -
//schematic
// LAST TIME SAVED: Jul 16 18:10:58 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module ice1f_array_RGT_IO_top12io ( cf_r, fabric_out_09, fabric_out_10,
     fabric_out_11, fabric_out_12, fabric_out_13, fabric_out_14,
     fabric_out_15, fabric_out_16, padeb, pado, sdo, slf_op_13_09,
     slf_op_13_10, slf_op_13_11, slf_op_13_12, slf_op_13_13,
     slf_op_13_14, slf_op_13_15, slf_op_13_16, spi_ss_in_b,
     SP4_h_l_13_09, SP4_h_l_13_10, SP4_h_l_13_11, SP4_h_l_13_12,
     SP4_h_l_13_13, SP4_h_l_13_14, SP4_h_l_13_15, SP4_h_l_13_16,
     SP12_h_l_13_09, SP12_h_l_13_10, SP12_h_l_13_11, SP12_h_l_13_12,
     SP12_h_l_13_13, SP12_h_l_13_14, SP12_h_l_13_15, SP12_h_l_13_16,
     bl, pgate, reset_b, sp4_v_b_13_09, sp4_v_t_41_40, vdd_cntl, wl,
     bnl_op_13_09, bs_en, cdone_in, ceb, glb_netwk_col, hiz_b, hold,
     lft_op_13_09, lft_op_13_10, lft_op_13_11, lft_op_13_12,
     lft_op_13_13, lft_op_13_14, lft_op_13_15, lft_op_13_16, mode,
     padin, prog, r, sdi, shift, spioeb, spiout, tclk, tnl_op_41_40,
     update );
output  fabric_out_09, fabric_out_10, fabric_out_11, fabric_out_12,
     fabric_out_13, fabric_out_14, fabric_out_15, fabric_out_16, sdo;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_13_12;
output [3:0]  slf_op_13_15;
output [3:0]  slf_op_13_14;
output [3:0]  slf_op_13_13;
output [3:0]  slf_op_13_16;
output [3:0]  slf_op_13_11;
output [3:0]  slf_op_13_10;
output [191:0]  cf_r;
output [11:0]  padeb;
output [11:0]  pado;
output [15:0]  spi_ss_in_b;
output [3:0]  slf_op_13_09;

inout [17:0]  bl;
inout [47:0]  SP4_h_l_13_09;
inout [47:0]  SP4_h_l_13_13;
inout [23:0]  SP12_h_l_13_13;
inout [47:0]  SP4_h_l_13_12;
inout [47:0]  SP4_h_l_13_15;
inout [47:0]  SP4_h_l_13_10;
inout [23:0]  SP12_h_l_13_09;
inout [15:0]  sp4_v_b_13_09;
inout [23:0]  SP12_h_l_13_11;
inout [23:0]  SP12_h_l_13_10;
inout [23:0]  SP12_h_l_13_15;
inout [23:0]  SP12_h_l_13_14;
inout [47:0]  SP4_h_l_13_14;
inout [23:0]  SP12_h_l_13_12;
inout [127:0]  pgate;
inout [23:0]  SP12_h_l_13_16;
inout [127:0]  vdd_cntl;
inout [127:0]  reset_b;
inout [15:0]  sp4_v_t_41_40;
inout [47:0]  SP4_h_l_13_11;
inout [127:0]  wl;
inout [47:0]  SP4_h_l_13_16;

input [7:0]  tnl_op_41_40;
input [7:0]  lft_op_13_15;
input [7:0]  lft_op_13_12;
input [7:0]  lft_op_13_14;
input [7:0]  lft_op_13_10;
input [7:0]  bnl_op_13_09;
input [7:0]  lft_op_13_09;
input [7:0]  lft_op_13_16;
input [7:0]  glb_netwk_col;
input [15:0]  spioeb;
input [11:0]  padin;
input [7:0]  lft_op_13_11;
input [16:9]  cdone_in;
input [7:0]  lft_op_13_13;
input [15:0]  spiout;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net625;

wire  [0:1]  net486;

wire  [0:15]  net416;

wire  [0:15]  net452;

wire  [7:0]  colbuf_cntl_b;

wire  [0:15]  net380;

wire  [0:15]  net524;

wire  [0:15]  net596;

wire  [7:0]  glb_netwk_t;

wire  [0:7]  net624;

wire  [7:0]  colbuf_cntl_t;

wire  [0:15]  net488;

wire  [0:7]  net626;

wire  [0:7]  net627;

wire  [0:7]  net629;

wire  [0:1]  net343;

wire  [0:15]  net560;

wire  [0:1]  net487;

wire  [0:7]  net628;

wire  [0:1]  net342;

wire  [7:0]  glb_netwk_b;



io_col4_RGT_rev I_io_13_16 ( .cbit_colcntl(net626[0:7]), .ceb(ceb),
     .sdo(sdo), .sdi(net365), .spiout(spiout[15:14]),
     .cdone_in(cdone_in[16]), .spioeb(spioeb[15:14]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(net342[0:1]), .pado(net342[0:1]),
     .padeb(net343[0:1]), .sp4_v_t(sp4_v_t_41_40[15:0]),
     .sp4_h_l(SP4_h_l_13_16[47:0]), .sp12_h_l(SP12_h_l_13_16[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[15:14]),
     .tnl_op(tnl_op_41_40[7:0]), .lft_op(lft_op_13_16[7:0]),
     .bnl_op(lft_op_13_15[7:0]), .pgate(pgate[127:112]),
     .reset(reset_b[127:112]), .sp4_v_b(net380[0:15]),
     .wl(wl[127:112]), .cf(cf_r[191:168]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[127:112]), .slf_op(slf_op_13_16[3:0]),
     .glb_netwk(glb_netwk_t[7:0]), .hold(hold),
     .fabric_out(fabric_out_16));
io_col4_RGT_rev I_io_13_15 ( .cbit_colcntl(net628[0:7]), .ceb(ceb),
     .sdo(net365), .sdi(net437), .spiout(spiout[13:12]),
     .cdone_in(cdone_in[15]), .spioeb(spioeb[13:12]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[11:10]), .pado(pado[11:10]),
     .padeb(padeb[11:10]), .sp4_v_t(net380[0:15]),
     .sp4_h_l(SP4_h_l_13_15[47:0]), .sp12_h_l(SP12_h_l_13_15[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[13:12]),
     .tnl_op(lft_op_13_16[7:0]), .lft_op(lft_op_13_15[7:0]),
     .bnl_op(lft_op_13_14[7:0]), .pgate(pgate[111:96]),
     .reset(reset_b[111:96]), .sp4_v_b(net452[0:15]), .wl(wl[111:96]),
     .cf(cf_r[167:144]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_13_15[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_15));
io_col4_RGT_rev I_io_13_13 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net401), .sdi(net581), .spiout(spiout[9:8]),
     .cdone_in(cdone_in[13]), .spioeb(spioeb[9:8]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[7:6]), .pado(pado[7:6]),
     .padeb(padeb[7:6]), .sp4_v_t(net416[0:15]),
     .sp4_h_l(SP4_h_l_13_13[47:0]), .sp12_h_l(SP12_h_l_13_13[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[9:8]),
     .tnl_op(lft_op_13_14[7:0]), .lft_op(lft_op_13_13[7:0]),
     .bnl_op(lft_op_13_12[7:0]), .pgate(pgate[79:64]),
     .reset(reset_b[79:64]), .sp4_v_b(net596[0:15]), .wl(wl[79:64]),
     .cf(cf_r[119:96]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_13_13[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_13));
io_col4_RGT_rev I_io_13_14 ( .cbit_colcntl(net627[0:7]), .ceb(ceb),
     .sdo(net437), .sdi(net401), .spiout(spiout[11:10]),
     .cdone_in(cdone_in[14]), .spioeb(spioeb[11:10]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[9:8]), .pado(pado[9:8]),
     .padeb(padeb[9:8]), .sp4_v_t(net452[0:15]),
     .sp4_h_l(SP4_h_l_13_14[47:0]), .sp12_h_l(SP12_h_l_13_14[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[11:10]),
     .tnl_op(lft_op_13_15[7:0]), .lft_op(lft_op_13_14[7:0]),
     .bnl_op(lft_op_13_13[7:0]), .pgate(pgate[95:80]),
     .reset(reset_b[95:80]), .sp4_v_b(net416[0:15]), .wl(wl[95:80]),
     .cf(cf_r[143:120]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_13_14[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_14));
io_col4_RGT_rev I_io_13_10 ( .cbit_colcntl(net624[0:7]), .ceb(ceb),
     .sdo(net473), .sdi(net509), .spiout(spiout[3:2]),
     .cdone_in(cdone_in[10]), .spioeb(spioeb[3:2]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(net486[0:1]), .pado(net486[0:1]),
     .padeb(net487[0:1]), .sp4_v_t(net488[0:15]),
     .sp4_h_l(SP4_h_l_13_10[47:0]), .sp12_h_l(SP12_h_l_13_10[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[3:2]),
     .tnl_op(lft_op_13_11[7:0]), .lft_op(lft_op_13_10[7:0]),
     .bnl_op(lft_op_13_09[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b(net524[0:15]), .wl(wl[31:16]),
     .cf(cf_r[47:24]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_13_10[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_10));
io_col4_RGT_rev I_io_13_09 ( .cbit_colcntl(net629[0:7]), .ceb(ceb),
     .sdo(net509), .sdi(sdi), .spiout(spiout[1:0]),
     .cdone_in(cdone_in[9]), .spioeb(spioeb[1:0]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .sp4_v_t(net524[0:15]),
     .sp4_h_l(SP4_h_l_13_09[47:0]), .sp12_h_l(SP12_h_l_13_09[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[1:0]),
     .tnl_op(lft_op_13_10[7:0]), .lft_op(lft_op_13_09[7:0]),
     .bnl_op(bnl_op_13_09[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(sp4_v_b_13_09[15:0]),
     .wl(wl[15:0]), .cf(cf_r[23:0]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_13_09[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold),
     .fabric_out(fabric_out_09));
io_col4_RGT_rev I_io_13_11 ( .cbit_colcntl(net625[0:7]), .ceb(ceb),
     .sdo(net545), .sdi(net473), .spiout(spiout[5:4]),
     .cdone_in(cdone_in[11]), .spioeb(spioeb[5:4]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[3:2]), .pado(pado[3:2]),
     .padeb(padeb[3:2]), .sp4_v_t(net560[0:15]),
     .sp4_h_l(SP4_h_l_13_11[47:0]), .sp12_h_l(SP12_h_l_13_11[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[5:4]),
     .tnl_op(lft_op_13_12[7:0]), .lft_op(lft_op_13_11[7:0]),
     .bnl_op(lft_op_13_10[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b(net488[0:15]), .wl(wl[47:32]),
     .cf(cf_r[71:48]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_13_11[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_11));
io_col4_RGT_rev I_io_13_12 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net581), .sdi(net545), .spiout(spiout[7:6]),
     .cdone_in(cdone_in[12]), .spioeb(spioeb[7:6]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[5:4]), .pado(pado[5:4]),
     .padeb(padeb[5:4]), .sp4_v_t(net596[0:15]),
     .sp4_h_l(SP4_h_l_13_12[47:0]), .sp12_h_l(SP12_h_l_13_12[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[7:6]),
     .tnl_op(lft_op_13_13[7:0]), .lft_op(lft_op_13_12[7:0]),
     .bnl_op(lft_op_13_11[7:0]), .pgate(pgate[63:48]),
     .reset(reset_b[63:48]), .sp4_v_b(net560[0:15]), .wl(wl[63:48]),
     .cf(cf_r[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_13_12[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_12));
clk_colbuf1kx8 I_clk_colbuf1kx8b ( .colbuf_cntl(colbuf_cntl_b[7:0]),
     .col_clk(glb_netwk_b[7:0]), .clk_in(glb_netwk_col[7:0]));
clk_colbuf1kx8 I_clk_colbuf1kx8t ( .colbuf_cntl(colbuf_cntl_t[7:0]),
     .col_clk(glb_netwk_t[7:0]), .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - io, Cell - io_col4_TOP_rev, View - schematic
// LAST TIME SAVED: Jul 10 10:35:31 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module io_col4_TOP_rev ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [23:0]  cf;
output [1:0]  spi_ss_in_b;
output [3:0]  slf_op;
output [1:0]  padeb;

inout [15:0]  sp4_v_t;
inout [17:0]  bl;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;

input [1:0]  padin;
input [1:0]  spioeb;
input [15:0]  wl;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [7:0]  glb_netwk;
input [1:0]  spiout;
input [15:0]  reset;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [0:7]  net0138;



ioe_col2rev I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .dout(slf_op[3:0]), .outclk(outclk), .hold(hold),
     .rstio(r), .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]}), .reset({reset[14], reset[15], reset[12], reset[13],
     reset[10], reset[11], reset[8], reset[9], reset[6], reset[7],
     reset[4], reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net128), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));
sbox1_colbdlc_rev Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net128));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net128));
rm6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net128, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .cbit_colcntl(net0138[0:7]),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min7({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}), .min5({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14], wl[15],
     wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4],
     wl[5], wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .prog(net128),
     .lc_trk_g1(lc_trk_g1[7:0]));

endmodule
// Library - leafcell, Cell - ice1f_array_TOP_IO_rgt, View - schematic
// LAST TIME SAVED: Jun 30 15:01:35 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module ice1f_array_TOP_IO_rgt ( bs_en_o, ceb_o, cf_top_l,
     fabric_out_07_17, fabric_out_08_17, hiz_b_o, mode_o, padeb_t_r,
     pado_t_r, r_o, sdo, shift_o, slf_op_07_17, slf_op_08_17,
     slf_op_09_17, slf_op_10_17, slf_op_11_17, slf_op_12_17, tclk_o,
     update_o, bl_07, bl_08, bl_09, bl_10, bl_11, bl_12, sp4_h_l_07_17,
     sp4_h_r_12_17, sp4_v_b_07_17, sp4_v_b_08_17, sp4_v_b_09_17,
     sp4_v_b_10_17, sp4_v_b_11_17, sp4_v_b_12_17, sp12_v_b_07_17,
     sp12_v_b_08_17, sp12_v_b_09_17, sp12_v_b_10_17, sp12_v_b_11_17,
     sp12_v_b_12_17, bnl_op_07_17, bnr_op_12_17, bs_en_i, ceb_i,
     end_of_startup_top_l, glb_net_07, glb_net_08, glb_net_09,
     glb_net_10, glb_net_11, glb_net_12, hiz_b_i, hold_t_r,
     lft_op_07_17, lft_op_08_17, lft_op_09_17, lft_op_10_17,
     lft_op_11_17, lft_op_12_17, mode_i, padin_t_r, pgate_l, prog, r_i,
     reset_l, sdi, shift_i, tclk_i, tiegnd, tievdd, update_i,
     vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_07_17, fabric_out_08_17, hiz_b_o,
     mode_o, r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_r, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, tiegnd, tievdd, update_i;

output [3:0]  slf_op_09_17;
output [3:0]  slf_op_11_17;
output [3:0]  slf_op_07_17;
output [3:0]  slf_op_12_17;
output [3:0]  slf_op_10_17;
output [3:0]  slf_op_08_17;
output [11:0]  padeb_t_r;
output [11:0]  pado_t_r;
output [143:0]  cf_top_l;

inout [15:0]  sp4_h_r_12_17;
inout [23:0]  sp12_v_b_10_17;
inout [23:0]  sp12_v_b_11_17;
inout [47:0]  sp4_v_b_11_17;
inout [47:0]  sp4_v_b_12_17;
inout [47:0]  sp4_v_b_09_17;
inout [47:0]  sp4_v_b_10_17;
inout [23:0]  sp12_v_b_07_17;
inout [47:0]  sp4_v_b_08_17;
inout [15:0]  sp4_h_l_07_17;
inout [23:0]  sp12_v_b_08_17;
inout [47:0]  sp4_v_b_07_17;
inout [23:0]  sp12_v_b_09_17;
inout [53:0]  bl_12;
inout [23:0]  sp12_v_b_12_17;
inout [53:0]  bl_08;
inout [53:0]  bl_09;
inout [53:0]  bl_07;
inout [41:0]  bl_10;
inout [53:0]  bl_11;

input [7:0]  lft_op_09_17;
input [7:0]  lft_op_11_17;
input [7:0]  glb_net_09;
input [7:0]  glb_net_11;
input [7:0]  lft_op_12_17;
input [15:0]  reset_l;
input [7:0]  lft_op_10_17;
input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_08;
input [7:0]  bnl_op_07_17;
input [15:0]  wl_l;
input [7:0]  glb_net_10;
input [7:0]  glb_net_07;
input [11:0]  padin_t_r;
input [7:0]  bnr_op_12_17;
input [7:0]  glb_net_12;
input [7:0]  lft_op_07_17;
input [7:0]  lft_op_08_17;
input [15:0]  pgate_l;
input [6:1]  end_of_startup_top_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net321;

wire  [0:15]  net317;

wire  [0:15]  net352;

wire  [0:1]  net503;

wire  [0:1]  net510;

wire  [0:15]  net387;

wire  [0:1]  net507;

wire  [0:15]  net282;

wire  [0:1]  net499;

wire  [0:15]  net422;

wire  [0:1]  net426;



io_col4_TOP_rev I_io_t07 ( .sdo(net479), .sdi(net267), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[1]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_07_17[15:0]), .mode(mode_i),
     .shift(shift_i), .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i),
     .tclk(tclk_i), .update(update_i), .padin(padin_t_r[1:0]),
     .pado(pado_t_r[1:0]), .padeb(padeb_t_r[1:0]),
     .sp4_v_b(net282[0:15]), .sp4_h_l(sp4_v_b_07_17[47:0]),
     .sp12_h_l(sp12_v_b_07_17[23:0]), .prog(prog),
     .spi_ss_in_b(net507[0:1]), .tnl_op(bnl_op_07_17[7:0]),
     .lft_op(lft_op_07_17[7:0]), .bnl_op(lft_op_08_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_07[5],
     bl_07[4], bl_07[37], bl_07[36], bl_07[35], bl_07[34], bl_07[33],
     bl_07[32], bl_07[14], bl_07[20], bl_07[19], bl_07[18], bl_07[17],
     bl_07[16], bl_07[27], bl_07[26], bl_07[25], bl_07[23]}),
     .wl(wl_l[15:0]), .cf(cf_top_l[23:0]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_07_17[3:0]),
     .glb_netwk(glb_net_07[7:0]), .hold(hold_t_r),
     .fabric_out(fabric_out_07_17));
io_col4_TOP_rev I_io_t08 ( .sdo(net267), .sdi(net302), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[2]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net282[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_r[3:2]), .pado(pado_t_r[3:2]),
     .padeb(padeb_t_r[3:2]), .sp4_v_b(net317[0:15]),
     .sp4_h_l(sp4_v_b_08_17[47:0]), .sp12_h_l(sp12_v_b_08_17[23:0]),
     .prog(prog), .spi_ss_in_b(net321[0:1]),
     .tnl_op(lft_op_07_17[7:0]), .lft_op(lft_op_08_17[7:0]),
     .bnl_op(lft_op_09_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_08[5], bl_08[4], bl_08[37],
     bl_08[36], bl_08[35], bl_08[34], bl_08[33], bl_08[32], bl_08[14],
     bl_08[20], bl_08[19], bl_08[18], bl_08[17], bl_08[16], bl_08[27],
     bl_08[26], bl_08[25], bl_08[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[47:24]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_08_17[3:0]), .glb_netwk(glb_net_08[7:0]),
     .hold(hold_t_r), .fabric_out(fabric_out_08_17));
io_col4_TOP_rev I_io_t09 ( .sdo(net302), .sdi(net337), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[3]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net317[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_r[5:4]), .pado(pado_t_r[5:4]),
     .padeb(padeb_t_r[5:4]), .sp4_v_b(net352[0:15]),
     .sp4_h_l(sp4_v_b_09_17[47:0]), .sp12_h_l(sp12_v_b_09_17[23:0]),
     .prog(prog), .spi_ss_in_b(net499[0:1]),
     .tnl_op(lft_op_08_17[7:0]), .lft_op(lft_op_09_17[7:0]),
     .bnl_op(lft_op_10_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_09[5], bl_09[4], bl_09[37],
     bl_09[36], bl_09[35], bl_09[34], bl_09[33], bl_09[32], bl_09[14],
     bl_09[20], bl_09[19], bl_09[18], bl_09[17], bl_09[16], bl_09[27],
     bl_09[26], bl_09[25], bl_09[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[71:48]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_09_17[3:0]), .glb_netwk(glb_net_09[7:0]),
     .hold(hold_t_r), .fabric_out(net370));
io_col4_TOP_rev I_io_t11 ( .sdo(net407), .sdi(net372), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[5]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net422[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_r[9:8]), .pado(pado_t_r[9:8]),
     .padeb(padeb_t_r[9:8]), .sp4_v_b(net387[0:15]),
     .sp4_h_l(sp4_v_b_11_17[47:0]), .sp12_h_l(sp12_v_b_11_17[23:0]),
     .prog(prog), .spi_ss_in_b(net503[0:1]),
     .tnl_op(lft_op_10_17[7:0]), .lft_op(lft_op_11_17[7:0]),
     .bnl_op(lft_op_12_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_11[5], bl_11[4], bl_11[37],
     bl_11[36], bl_11[35], bl_11[34], bl_11[33], bl_11[32], bl_11[14],
     bl_11[20], bl_11[19], bl_11[18], bl_11[17], bl_11[16], bl_11[27],
     bl_11[26], bl_11[25], bl_11[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[119:96]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_11_17[3:0]), .glb_netwk(glb_net_11[7:0]),
     .hold(hold_t_r), .fabric_out(net405));
io_col4_TOP_rev I_io_t10 ( .sdo(net337), .sdi(net407), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[4]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net352[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_r[7:6]), .pado(pado_t_r[7:6]),
     .padeb(padeb_t_r[7:6]), .sp4_v_b(net422[0:15]),
     .sp4_h_l(sp4_v_b_10_17[47:0]), .sp12_h_l(sp12_v_b_10_17[23:0]),
     .prog(prog), .spi_ss_in_b(net426[0:1]),
     .tnl_op(lft_op_09_17[7:0]), .lft_op(lft_op_10_17[7:0]),
     .bnl_op(lft_op_11_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_10[5], bl_10[4], bl_10[37],
     bl_10[36], bl_10[35], bl_10[34], bl_10[33], bl_10[32], bl_10[14],
     bl_10[20], bl_10[19], bl_10[18], bl_10[17], bl_10[16], bl_10[27],
     bl_10[26], bl_10[25], bl_10[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[95:72]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_10_17[3:0]), .glb_netwk(glb_net_10[7:0]),
     .hold(hold_t_r), .fabric_out(net440));
io_col4_TOP_rev I_io_t12 ( .sdo(net372), .sdi(sdi), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[6]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net387[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_r[11:10]),
     .pado(pado_t_r[11:10]), .padeb(padeb_t_r[11:10]),
     .sp4_v_b(sp4_h_r_12_17[15:0]), .sp4_h_l(sp4_v_b_12_17[47:0]),
     .sp12_h_l(sp12_v_b_12_17[23:0]), .prog(prog),
     .spi_ss_in_b(net510[0:1]), .tnl_op(lft_op_11_17[7:0]),
     .lft_op(lft_op_12_17[7:0]), .bnl_op(bnr_op_12_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_12[5],
     bl_12[4], bl_12[37], bl_12[36], bl_12[35], bl_12[34], bl_12[33],
     bl_12[32], bl_12[14], bl_12[20], bl_12[19], bl_12[18], bl_12[17],
     bl_12[16], bl_12[27], bl_12[26], bl_12[25], bl_12[23]}),
     .wl(wl_l[15:0]), .cf(cf_top_l[143:120]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_12_17[3:0]),
     .glb_netwk(glb_net_12[7:0]), .hold(hold_t_r),
     .fabric_out(net509));
scanbuf1f I_scanbuf_mt ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(net479), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(tclk_o), .shift_o(shift_o),
     .sdo(sdo), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));

endmodule
// Library - leafcell, Cell - bram_4k_sr_bankin, View - schematic
// LAST TIME SAVED: Aug 15 18:05:22 2007
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module bram_4k_sr_bankin ( bm_dm, bm_sweb, clk, rcapmux_en, rst, bm_q,
     bm_sdi, wdummymux_en );

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(net150), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));
ml_mux2_hvt_schematic I20 ( .in1(wdummy_reg), .in0(bm_dm[0]),
     .out(net150), .sel(wdummymux_en));
leafcell_ml_dff_schematic I19 ( .R(rst), .D(bm_sdi), .CLK(clk),
     .QN(net157), .Q(wdummy_reg));

endmodule
// Library - leafcell, Cell - bram_4k_bankin, View - schematic
// LAST TIME SAVED: Aug 15 18:08:05 2007
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module bram_4k_bankin ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_ab;
input [7:0]  bm_sa;
input [7:0]  bm_aa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [14:0]  bm_dm;



tielo I15 ( .tielo(net102));
tielo I18 ( .tielo(net103));
bram_4k_sr_bankin I12 ( .bm_dm({bm_sdo, bm_dm[14:0]}), .rst(net103),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM({bm_sdo, bm_dm[14:0]}), .WEBM(bm_sweb), .WEB(web),
     .REBM(bm_sreb), .REB(reb), .D(bm_d[15:0]), .CLKW(net82),
     .CLKR(net80), .BWEBM({net102, net102, net102, net102, net102,
     net102, net102, net102, net102, net102, net102, net102, net102,
     net102, net102, net102}), .BWEB(bm_bweb[15:0]), .BIST(bm_init),
     .AMB(bm_sa[7:0]), .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]),
     .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net98), .out(net80));
bram_bufferx6 I8 ( .in(net94), .out(net82));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net94), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net98), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - leafcell, Cell - bram_4kbankin_pbuffer_top, View -
//schematic
// LAST TIME SAVED: Aug 24 17:33:59 2007
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module bram_4kbankin_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [7:0]  bm_sa_o;
output [15:0]  bm_q;

input [7:0]  bm_sa_i;
input [7:0]  bm_ab;
input [7:0]  bm_aa;
input [15:0]  bm_d;
input [15:0]  bm_bweb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k_bankin I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - leafcell, Cell - bram_4kprouting_tbankin, View - schematic
// LAST TIME SAVED: Jan  8 10:39:02 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module bram_4kprouting_tbankin ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;

inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_v_t_top;
inout [23:0]  sp12_h_l_top;
inout [23:0]  sp12_v_t_top;
inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [41:0]  bl;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_v_b_top;

input [7:0]  glb_netwk;
input [7:0]  tnr_op_bot;
input [7:0]  rgt_op_top;
input [7:0]  bnl_op_bot;
input [7:0]  lft_op_bot;
input [7:0]  tnl_op_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  lft_op_top;
input [7:0]  tnr_op_top;
input [15:0]  pgate_bot;
input [7:0]  bnl_op_top;
input [7:0]  top_op_top;
input [7:0]  bot_op_bot;
input [15:0]  vdd_cntl_top;
input [7:0]  bnr_op_bot;
input [7:0]  bnr_op_top;
input [15:0]  reset_b_top;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_bot;
input [15:0]  wl_top;
input [15:0]  wl_bot;
input [15:0]  pgate_top;
input [7:0]  rgt_op_bot;
input [15:0]  reset_b_bot;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net210;

wire  [0:7]  net316;

wire  [0:7]  net208;

wire  [0:7]  net295;

wire  [0:7]  net211;

wire  [7:0]  in2_top;

wire  [0:7]  net242;

wire  [0:7]  net209;

wire  [0:7]  net243;

wire  [0:7]  net0240;

wire  [0:7]  net0208;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net240;

wire  [15:0]  bm_bweb;

wire  [0:7]  net241;

wire  [7:0]  in2_bot;

wire  [15:0]  bm_d;



bram_routing_tracks4rev12 I_bot ( .cbit_colcntl(net0208[0:7]),
     .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15], vdd_cntl_bot[12],
     vdd_cntl_bot[13], vdd_cntl_bot[10], vdd_cntl_bot[11],
     vdd_cntl_bot[8], vdd_cntl_bot[9], vdd_cntl_bot[6],
     vdd_cntl_bot[7], vdd_cntl_bot[4], vdd_cntl_bot[5],
     vdd_cntl_bot[2], vdd_cntl_bot[3], vdd_cntl_bot[0],
     vdd_cntl_bot[1]}), .s_r(net213), .wl({wl_bot[14], wl_bot[15],
     wl_bot[12], wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8],
     wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2],
     wl_bot[3], wl_bot[0], wl_bot[1]}), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev12 I_top ( .cbit_colcntl(net0240[0:7]),
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .s_r(net245), .wl({wl_top[14], wl_top[15],
     wl_top[12], wl_top[13], wl_top[10], wl_top[11], wl_top[8],
     wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2],
     wl_top[3], wl_top[0], wl_top[1]}), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbankin_pbuffer_top I_bram_4kbankin_pbuffer_top (
     .bm_q({slf_op_top[7:0], slf_op_bot[7:0]}),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_init_i(bm_init_i),
     .bm_ren(net245), .bm_wen(net213), .bm_d(bm_d[15:0]),
     .bm_clkr(net244), .bm_clkw(net212), .bm_bweb(bm_bweb[15:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sdo_o(bm_sdo_o),
     .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sdo_i(bm_sdo_i), .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i),
     .bm_sdi_o(bm_sdi_o), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_aa(net295[0:7]), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_sweb_o(bm_sweb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_b ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}),
     .bl(bl[41:26]), .wl({wl_bot[14], wl_bot[15], wl_bot[12],
     wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8], wl_bot[9],
     wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2], wl_bot[3],
     wl_bot[0], wl_bot[1]}), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .op(slf_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .sp12_h_r({sp12_h_r_bot[22],
     sp12_h_r_bot[6], sp12_h_r_bot[20], sp12_h_r_bot[4],
     sp12_h_r_bot[18], sp12_h_r_bot[2], sp12_h_r_bot[16],
     sp12_h_r_bot[0], sp12_h_r_bot[14], sp12_h_r_bot[12],
     sp12_h_r_bot[10], sp12_h_r_bot[8]}), .sp4_v_b({sp4_v_b_bot[46],
     sp4_v_b_bot[30], sp4_v_b_bot[14], sp4_v_b_bot[44],
     sp4_v_b_bot[28], sp4_v_b_bot[12], sp4_v_b_bot[42],
     sp4_v_b_bot[26], sp4_v_b_bot[10], sp4_v_b_bot[40],
     sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38], sp4_v_b_bot[22],
     sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20], sp4_v_b_bot[4],
     sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2], sp4_v_b_bot[32],
     sp4_v_b_bot[16], sp4_v_b_bot[0]}), .sp4_r_v_b({sp4_r_v_b_bot[47],
     sp4_r_v_b_bot[31], sp4_r_v_b_bot[15], sp4_r_v_b_bot[45],
     sp4_r_v_b_bot[29], sp4_r_v_b_bot[13], sp4_r_v_b_bot[43],
     sp4_r_v_b_bot[27], sp4_r_v_b_bot[11], sp4_r_v_b_bot[41],
     sp4_r_v_b_bot[25], sp4_r_v_b_bot[9], sp4_r_v_b_bot[39],
     sp4_r_v_b_bot[23], sp4_r_v_b_bot[7], sp4_r_v_b_bot[37],
     sp4_r_v_b_bot[21], sp4_r_v_b_bot[5], sp4_r_v_b_bot[35],
     sp4_r_v_b_bot[19], sp4_r_v_b_bot[3], sp4_r_v_b_bot[33],
     sp4_r_v_b_bot[17], sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46],
     sp4_h_r_bot[30], sp4_h_r_bot[14], sp4_h_r_bot[44],
     sp4_h_r_bot[28], sp4_h_r_bot[12], sp4_h_r_bot[42],
     sp4_h_r_bot[26], sp4_h_r_bot[10], sp4_h_r_bot[40],
     sp4_h_r_bot[24], sp4_h_r_bot[8], sp4_h_r_bot[38], sp4_h_r_bot[22],
     sp4_h_r_bot[6], sp4_h_r_bot[36], sp4_h_r_bot[20], sp4_h_r_bot[4],
     sp4_h_r_bot[34], sp4_h_r_bot[18], sp4_h_r_bot[2], sp4_h_r_bot[32],
     sp4_h_r_bot[16], sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]),
     .in2(in2_bot[7:0]), .in1(bm_d[7:0]), .in0(net295[0:7]),
     .sp12_v_b({sp12_v_b_bot[14], sp12_v_b_bot[12], sp12_v_b_bot[10],
     sp12_v_b_bot[8], sp12_v_b_bot[22], sp12_v_b_bot[6],
     sp12_v_b_bot[20], sp12_v_b_bot[4], sp12_v_b_bot[18],
     sp12_v_b_bot[2], sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_t ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}),
     .bl(bl[41:26]), .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12],
     sp12_v_b_top[10], sp12_v_b_top[8], sp12_v_b_top[22],
     sp12_v_b_top[6], sp12_v_b_top[20], sp12_v_b_top[4],
     sp12_v_b_top[18], sp12_v_b_top[2], sp12_v_b_top[16],
     sp12_v_b_top[0]}), .wl({wl_top[14], wl_top[15], wl_top[12],
     wl_top[13], wl_top[10], wl_top[11], wl_top[8], wl_top[9],
     wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2], wl_top[3],
     wl_top[0], wl_top[1]}), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .op(slf_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .sp12_h_r({sp12_h_r_top[22],
     sp12_h_r_top[6], sp12_h_r_top[20], sp12_h_r_top[4],
     sp12_h_r_top[18], sp12_h_r_top[2], sp12_h_r_top[16],
     sp12_h_r_top[0], sp12_h_r_top[14], sp12_h_r_top[12],
     sp12_h_r_top[10], sp12_h_r_top[8]}), .sp4_v_b({sp4_v_b_top[46],
     sp4_v_b_top[30], sp4_v_b_top[14], sp4_v_b_top[44],
     sp4_v_b_top[28], sp4_v_b_top[12], sp4_v_b_top[42],
     sp4_v_b_top[26], sp4_v_b_top[10], sp4_v_b_top[40],
     sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38], sp4_v_b_top[22],
     sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20], sp4_v_b_top[4],
     sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2], sp4_v_b_top[32],
     sp4_v_b_top[16], sp4_v_b_top[0]}), .sp4_r_v_b({sp4_r_v_b_top[47],
     sp4_r_v_b_top[31], sp4_r_v_b_top[15], sp4_r_v_b_top[45],
     sp4_r_v_b_top[29], sp4_r_v_b_top[13], sp4_r_v_b_top[43],
     sp4_r_v_b_top[27], sp4_r_v_b_top[11], sp4_r_v_b_top[41],
     sp4_r_v_b_top[25], sp4_r_v_b_top[9], sp4_r_v_b_top[39],
     sp4_r_v_b_top[23], sp4_r_v_b_top[7], sp4_r_v_b_top[37],
     sp4_r_v_b_top[21], sp4_r_v_b_top[5], sp4_r_v_b_top[35],
     sp4_r_v_b_top[19], sp4_r_v_b_top[3], sp4_r_v_b_top[33],
     sp4_r_v_b_top[17], sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46],
     sp4_h_r_top[30], sp4_h_r_top[14], sp4_h_r_top[44],
     sp4_h_r_top[28], sp4_h_r_top[12], sp4_h_r_top[42],
     sp4_h_r_top[26], sp4_h_r_top[10], sp4_h_r_top[40],
     sp4_h_r_top[24], sp4_h_r_top[8], sp4_h_r_top[38], sp4_h_r_top[22],
     sp4_h_r_top[6], sp4_h_r_top[36], sp4_h_r_top[20], sp4_h_r_top[4],
     sp4_h_r_top[34], sp4_h_r_top[18], sp4_h_r_top[2], sp4_h_r_top[32],
     sp4_h_r_top[16], sp4_h_r_top[0]}), .in3(bm_bweb[15:8]),
     .in2(in2_top[7:0]), .in1(bm_d[15:8]), .in0(net316[0:7]));

endmodule
// Library - leafcell, Cell - bram_4kbankout_pbuffer_top, View -
//schematic
// LAST TIME SAVED: Aug 24 17:34:59 2007
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module bram_4kbankout_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [7:0]  bm_sa_o;
output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_aa;
input [7:0]  bm_sa_i;
input [7:0]  bm_ab;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_4k_bankout I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));

endmodule
// Library - leafcell, Cell - bram_4kprouting_tbankout, View -
//schematic
// LAST TIME SAVED: Jan  8 10:42:36 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module bram_4kprouting_tbankout ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;

inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_h_l_top;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_r_v_b_bot;
inout [41:0]  bl;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_h_r_top;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_v_b_bot;

input [15:0]  pgate_top;
input [7:0]  bnr_op_top;
input [7:0]  bnl_op_bot;
input [15:0]  wl_bot;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_top;
input [7:0]  tnr_op_top;
input [7:0]  lft_op_bot;
input [7:0]  tnr_op_bot;
input [7:0]  rgt_op_top;
input [7:0]  bnr_op_bot;
input [7:0]  tnl_op_bot;
input [15:0]  reset_b_top;
input [15:0]  pgate_bot;
input [15:0]  reset_b_bot;
input [7:0]  lft_op_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  bnl_op_top;
input [7:0]  top_op_top;
input [7:0]  rgt_op_bot;
input [15:0]  vdd_cntl_top;
input [7:0]  glb_netwk;
input [7:0]  bot_op_bot;
input [15:0]  wl_top;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net208;

wire  [0:7]  net242;

wire  [0:7]  net240;

wire  [0:7]  net211;

wire  [0:7]  net243;

wire  [0:7]  net295;

wire  [0:7]  net241;

wire  [0:7]  net209;

wire  [0:7]  net0208;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net0240;

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [0:7]  net316;

wire  [15:0]  bm_d;

wire  [0:7]  net210;



bram_routing_tracks4rev12 I_bot ( .cbit_colcntl(net0208[0:7]),
     .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15], vdd_cntl_bot[12],
     vdd_cntl_bot[13], vdd_cntl_bot[10], vdd_cntl_bot[11],
     vdd_cntl_bot[8], vdd_cntl_bot[9], vdd_cntl_bot[6],
     vdd_cntl_bot[7], vdd_cntl_bot[4], vdd_cntl_bot[5],
     vdd_cntl_bot[2], vdd_cntl_bot[3], vdd_cntl_bot[0],
     vdd_cntl_bot[1]}), .s_r(net213), .wl({wl_bot[14], wl_bot[15],
     wl_bot[12], wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8],
     wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2],
     wl_bot[3], wl_bot[0], wl_bot[1]}), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev12 I_top ( .cbit_colcntl(net0240[0:7]),
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .s_r(net245), .wl({wl_top[14], wl_top[15],
     wl_top[12], wl_top[13], wl_top[10], wl_top[11], wl_top[8],
     wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2],
     wl_top[3], wl_top[0], wl_top[1]}), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbankout_pbuffer_top I_bram_4kbankout_pbuffer_top (
     .bm_q({slf_op_top[7:0], slf_op_bot[7:0]}),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_init_i(bm_init_i),
     .bm_ren(net245), .bm_wen(net213), .bm_d(bm_d[15:0]),
     .bm_clkr(net244), .bm_clkw(net212), .bm_bweb(bm_bweb[15:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sdo_o(bm_sdo_o),
     .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sdo_i(bm_sdo_i), .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i),
     .bm_sdi_o(bm_sdi_o), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_aa(net295[0:7]), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_sweb_o(bm_sweb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_b ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}),
     .bl(bl[41:26]), .wl({wl_bot[14], wl_bot[15], wl_bot[12],
     wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8], wl_bot[9],
     wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2], wl_bot[3],
     wl_bot[0], wl_bot[1]}), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .op(slf_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .sp12_h_r({sp12_h_r_bot[22],
     sp12_h_r_bot[6], sp12_h_r_bot[20], sp12_h_r_bot[4],
     sp12_h_r_bot[18], sp12_h_r_bot[2], sp12_h_r_bot[16],
     sp12_h_r_bot[0], sp12_h_r_bot[14], sp12_h_r_bot[12],
     sp12_h_r_bot[10], sp12_h_r_bot[8]}), .sp4_v_b({sp4_v_b_bot[46],
     sp4_v_b_bot[30], sp4_v_b_bot[14], sp4_v_b_bot[44],
     sp4_v_b_bot[28], sp4_v_b_bot[12], sp4_v_b_bot[42],
     sp4_v_b_bot[26], sp4_v_b_bot[10], sp4_v_b_bot[40],
     sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38], sp4_v_b_bot[22],
     sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20], sp4_v_b_bot[4],
     sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2], sp4_v_b_bot[32],
     sp4_v_b_bot[16], sp4_v_b_bot[0]}), .sp4_r_v_b({sp4_r_v_b_bot[47],
     sp4_r_v_b_bot[31], sp4_r_v_b_bot[15], sp4_r_v_b_bot[45],
     sp4_r_v_b_bot[29], sp4_r_v_b_bot[13], sp4_r_v_b_bot[43],
     sp4_r_v_b_bot[27], sp4_r_v_b_bot[11], sp4_r_v_b_bot[41],
     sp4_r_v_b_bot[25], sp4_r_v_b_bot[9], sp4_r_v_b_bot[39],
     sp4_r_v_b_bot[23], sp4_r_v_b_bot[7], sp4_r_v_b_bot[37],
     sp4_r_v_b_bot[21], sp4_r_v_b_bot[5], sp4_r_v_b_bot[35],
     sp4_r_v_b_bot[19], sp4_r_v_b_bot[3], sp4_r_v_b_bot[33],
     sp4_r_v_b_bot[17], sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46],
     sp4_h_r_bot[30], sp4_h_r_bot[14], sp4_h_r_bot[44],
     sp4_h_r_bot[28], sp4_h_r_bot[12], sp4_h_r_bot[42],
     sp4_h_r_bot[26], sp4_h_r_bot[10], sp4_h_r_bot[40],
     sp4_h_r_bot[24], sp4_h_r_bot[8], sp4_h_r_bot[38], sp4_h_r_bot[22],
     sp4_h_r_bot[6], sp4_h_r_bot[36], sp4_h_r_bot[20], sp4_h_r_bot[4],
     sp4_h_r_bot[34], sp4_h_r_bot[18], sp4_h_r_bot[2], sp4_h_r_bot[32],
     sp4_h_r_bot[16], sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]),
     .in2(in2_bot[7:0]), .in1(bm_d[7:0]), .in0(net295[0:7]),
     .sp12_v_b({sp12_v_b_bot[14], sp12_v_b_bot[12], sp12_v_b_bot[10],
     sp12_v_b_bot[8], sp12_v_b_bot[22], sp12_v_b_bot[6],
     sp12_v_b_bot[20], sp12_v_b_bot[4], sp12_v_b_bot[18],
     sp12_v_b_bot[2], sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_t ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}),
     .bl(bl[41:26]), .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12],
     sp12_v_b_top[10], sp12_v_b_top[8], sp12_v_b_top[22],
     sp12_v_b_top[6], sp12_v_b_top[20], sp12_v_b_top[4],
     sp12_v_b_top[18], sp12_v_b_top[2], sp12_v_b_top[16],
     sp12_v_b_top[0]}), .wl({wl_top[14], wl_top[15], wl_top[12],
     wl_top[13], wl_top[10], wl_top[11], wl_top[8], wl_top[9],
     wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2], wl_top[3],
     wl_top[0], wl_top[1]}), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .op(slf_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .sp12_h_r({sp12_h_r_top[22],
     sp12_h_r_top[6], sp12_h_r_top[20], sp12_h_r_top[4],
     sp12_h_r_top[18], sp12_h_r_top[2], sp12_h_r_top[16],
     sp12_h_r_top[0], sp12_h_r_top[14], sp12_h_r_top[12],
     sp12_h_r_top[10], sp12_h_r_top[8]}), .sp4_v_b({sp4_v_b_top[46],
     sp4_v_b_top[30], sp4_v_b_top[14], sp4_v_b_top[44],
     sp4_v_b_top[28], sp4_v_b_top[12], sp4_v_b_top[42],
     sp4_v_b_top[26], sp4_v_b_top[10], sp4_v_b_top[40],
     sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38], sp4_v_b_top[22],
     sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20], sp4_v_b_top[4],
     sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2], sp4_v_b_top[32],
     sp4_v_b_top[16], sp4_v_b_top[0]}), .sp4_r_v_b({sp4_r_v_b_top[47],
     sp4_r_v_b_top[31], sp4_r_v_b_top[15], sp4_r_v_b_top[45],
     sp4_r_v_b_top[29], sp4_r_v_b_top[13], sp4_r_v_b_top[43],
     sp4_r_v_b_top[27], sp4_r_v_b_top[11], sp4_r_v_b_top[41],
     sp4_r_v_b_top[25], sp4_r_v_b_top[9], sp4_r_v_b_top[39],
     sp4_r_v_b_top[23], sp4_r_v_b_top[7], sp4_r_v_b_top[37],
     sp4_r_v_b_top[21], sp4_r_v_b_top[5], sp4_r_v_b_top[35],
     sp4_r_v_b_top[19], sp4_r_v_b_top[3], sp4_r_v_b_top[33],
     sp4_r_v_b_top[17], sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46],
     sp4_h_r_top[30], sp4_h_r_top[14], sp4_h_r_top[44],
     sp4_h_r_top[28], sp4_h_r_top[12], sp4_h_r_top[42],
     sp4_h_r_top[26], sp4_h_r_top[10], sp4_h_r_top[40],
     sp4_h_r_top[24], sp4_h_r_top[8], sp4_h_r_top[38], sp4_h_r_top[22],
     sp4_h_r_top[6], sp4_h_r_top[36], sp4_h_r_top[20], sp4_h_r_top[4],
     sp4_h_r_top[34], sp4_h_r_top[18], sp4_h_r_top[2], sp4_h_r_top[32],
     sp4_h_r_top[16], sp4_h_r_top[0]}), .in3(bm_bweb[15:8]),
     .in2(in2_top[7:0]), .in1(bm_d[15:8]), .in0(net316[0:7]));

endmodule
// Library - leafcell, Cell - bram_4kbank_pbuffer_top, View - schematic
// LAST TIME SAVED: Aug 24 17:33:08 2007
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module bram_4kbank_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [7:0]  bm_sa_o;

input [15:0]  bm_bweb;
input [7:0]  bm_aa;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - misc, Cell - ml_osc_logic, View - schematic
// LAST TIME SAVED: Aug 28 08:48:45 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_osc_logic ( sel_trim, clkin, smc_osc_fsel, smc_oscen );

input  clkin, smc_oscen;

output [3:0]  sel_trim;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:2]  in_sel;



tiehi I280 ( .tiehi(net058));
ml_dff I174 ( .R(reset_ff), .D(net050), .CLK(clkin_buf_b), .QN(net150),
     .Q(net172));
ml_dff I238 ( .R(reset_ff), .D(net050), .CLK(clkin_buf), .QN(net154),
     .Q(net177));
ml_dff I244 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf),
     .QN(net155), .Q(net182));
ml_dff I245 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf_b),
     .QN(net153), .Q(net187));
ml_dff I242 ( .R(reset_ff), .D(net048), .CLK(clkin_buf_b), .QN(net191),
     .Q(net192));
ml_dff I243 ( .R(reset_ff), .D(net048), .CLK(clkin_buf), .QN(net152),
     .Q(net197));
ml_mux2_hvt I279 ( .in1(net182), .in0(net187), .out(sel_trim[0]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I277 ( .in1(net057), .in0(net061), .out(sel_trim[2]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I278 ( .in1(net052), .in0(net054), .out(sel_trim[1]),
     .sel(clkin_buf_delay));
nor2_hvt I256 ( .A(smc_osc_fsel[1]), .B(smc_osc_fsel[0]),
     .Y(in_sel[2]));
inv_hvt I263 ( .A(clkin_buf), .Y(net065));
inv_hvt I252 ( .A(smc_oscen), .Y(reset_ff));
inv_hvt I264 ( .A(net065), .Y(net063));
inv_hvt I253 ( .A(clkin_buf_b), .Y(clkin_buf));
inv_hvt I254 ( .A(clkin), .Y(clkin_buf_b));
inv_hvt I255 ( .A(smc_osc_fsel[1]), .Y(in_sel[1]));
inv_hvt I266 ( .A(net063), .Y(net059));
inv_hvt I265 ( .A(net059), .Y(net0143));
inv_hvt I274 ( .A(net177), .Y(net057));
inv_hvt I273 ( .A(net172), .Y(net061));
inv_hvt I275 ( .A(net192), .Y(net054));
inv_hvt I276 ( .A(net197), .Y(net052));
inv_hvt I261 ( .A(in_sel[2]), .Y(net050));
inv_hvt I267 ( .A(net0143), .Y(net0144));
inv_hvt I262 ( .A(in_sel[1]), .Y(net048));
inv_hvt I268 ( .A(net0144), .Y(net0145));
inv_hvt I269 ( .A(net0142), .Y(clkin_buf_delay));
inv_hvt I270 ( .A(net0145), .Y(net0142));
inv_hvt I176 ( .A(net058), .Y(sel_trim[3]));

endmodule
// Library - io, Cell - PVDD1DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:14:35 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module PVDD1DGZ ( VDD );
input  VDD;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - leafcell, Cell - bram_4kprouting_tbank, View - schematic
// LAST TIME SAVED: Jan  8 10:42:51 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module bram_4kprouting_tbank ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, cbit_colcntl, slf_op_bot, slf_op_top, bl,
     sp4_h_l_bot, sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  slf_op_top;
output [7:0]  slf_op_bot;
output [7:0]  cbit_colcntl;
output [7:0]  bm_sa_o;

inout [47:0]  sp4_v_t_top;
inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_h_l_bot;
inout [41:0]  bl;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_h_l_top;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_h_l_top;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_top;

input [7:0]  bnl_op_top;
input [7:0]  rgt_op_bot;
input [7:0]  tnr_op_bot;
input [7:0]  bot_op_bot;
input [7:0]  lft_op_bot;
input [7:0]  tnr_op_top;
input [7:0]  tnl_op_bot;
input [7:0]  top_op_top;
input [7:0]  glb_netwk;
input [7:0]  lft_op_top;
input [7:0]  bnl_op_bot;
input [15:0]  pgate_top;
input [15:0]  reset_b_bot;
input [15:0]  wl_bot;
input [15:0]  wl_top;
input [7:0]  bm_sa_i;
input [7:0]  rgt_op_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  bnr_op_top;
input [15:0]  pgate_bot;
input [15:0]  vdd_cntl_top;
input [7:0]  bnr_op_bot;
input [15:0]  reset_b_top;
input [7:0]  tnl_op_top;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net240;

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net209;

wire  [0:7]  net241;

wire  [0:7]  net211;

wire  [0:7]  net243;

wire  [0:7]  net316;

wire  [0:7]  net210;

wire  [0:7]  net208;

wire  [0:7]  net0240;

wire  [0:7]  net295;

wire  [0:7]  net242;



bram_routing_tracks4rev12 I_bot ( .cbit_colcntl(cbit_colcntl[7:0]),
     .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15], vdd_cntl_bot[12],
     vdd_cntl_bot[13], vdd_cntl_bot[10], vdd_cntl_bot[11],
     vdd_cntl_bot[8], vdd_cntl_bot[9], vdd_cntl_bot[6],
     vdd_cntl_bot[7], vdd_cntl_bot[4], vdd_cntl_bot[5],
     vdd_cntl_bot[2], vdd_cntl_bot[3], vdd_cntl_bot[0],
     vdd_cntl_bot[1]}), .s_r(net213), .wl({wl_bot[14], wl_bot[15],
     wl_bot[12], wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8],
     wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2],
     wl_bot[3], wl_bot[0], wl_bot[1]}), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev12 I_top ( .cbit_colcntl(net0240[0:7]),
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .s_r(net245), .wl({wl_top[14], wl_top[15],
     wl_top[12], wl_top[13], wl_top[10], wl_top[11], wl_top[8],
     wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2],
     wl_top[3], wl_top[0], wl_top[1]}), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbank_pbuffer_top I_bram_4kbank_pbuffer_top (
     .bm_q({slf_op_top[7:0], slf_op_bot[7:0]}),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_init_i(bm_init_i),
     .bm_ren(net245), .bm_wen(net213), .bm_d(bm_d[15:0]),
     .bm_clkr(net244), .bm_clkw(net212), .bm_bweb(bm_bweb[15:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sdo_o(bm_sdo_o),
     .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sdo_i(bm_sdo_i), .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i),
     .bm_sdi_o(bm_sdi_o), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_aa(net295[0:7]), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_sweb_o(bm_sweb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_b ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}),
     .bl(bl[41:26]), .wl({wl_bot[14], wl_bot[15], wl_bot[12],
     wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8], wl_bot[9],
     wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2], wl_bot[3],
     wl_bot[0], wl_bot[1]}), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .op(slf_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .sp12_h_r({sp12_h_r_bot[22],
     sp12_h_r_bot[6], sp12_h_r_bot[20], sp12_h_r_bot[4],
     sp12_h_r_bot[18], sp12_h_r_bot[2], sp12_h_r_bot[16],
     sp12_h_r_bot[0], sp12_h_r_bot[14], sp12_h_r_bot[12],
     sp12_h_r_bot[10], sp12_h_r_bot[8]}), .sp4_v_b({sp4_v_b_bot[46],
     sp4_v_b_bot[30], sp4_v_b_bot[14], sp4_v_b_bot[44],
     sp4_v_b_bot[28], sp4_v_b_bot[12], sp4_v_b_bot[42],
     sp4_v_b_bot[26], sp4_v_b_bot[10], sp4_v_b_bot[40],
     sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38], sp4_v_b_bot[22],
     sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20], sp4_v_b_bot[4],
     sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2], sp4_v_b_bot[32],
     sp4_v_b_bot[16], sp4_v_b_bot[0]}), .sp4_r_v_b({sp4_r_v_b_bot[47],
     sp4_r_v_b_bot[31], sp4_r_v_b_bot[15], sp4_r_v_b_bot[45],
     sp4_r_v_b_bot[29], sp4_r_v_b_bot[13], sp4_r_v_b_bot[43],
     sp4_r_v_b_bot[27], sp4_r_v_b_bot[11], sp4_r_v_b_bot[41],
     sp4_r_v_b_bot[25], sp4_r_v_b_bot[9], sp4_r_v_b_bot[39],
     sp4_r_v_b_bot[23], sp4_r_v_b_bot[7], sp4_r_v_b_bot[37],
     sp4_r_v_b_bot[21], sp4_r_v_b_bot[5], sp4_r_v_b_bot[35],
     sp4_r_v_b_bot[19], sp4_r_v_b_bot[3], sp4_r_v_b_bot[33],
     sp4_r_v_b_bot[17], sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46],
     sp4_h_r_bot[30], sp4_h_r_bot[14], sp4_h_r_bot[44],
     sp4_h_r_bot[28], sp4_h_r_bot[12], sp4_h_r_bot[42],
     sp4_h_r_bot[26], sp4_h_r_bot[10], sp4_h_r_bot[40],
     sp4_h_r_bot[24], sp4_h_r_bot[8], sp4_h_r_bot[38], sp4_h_r_bot[22],
     sp4_h_r_bot[6], sp4_h_r_bot[36], sp4_h_r_bot[20], sp4_h_r_bot[4],
     sp4_h_r_bot[34], sp4_h_r_bot[18], sp4_h_r_bot[2], sp4_h_r_bot[32],
     sp4_h_r_bot[16], sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]),
     .in2(in2_bot[7:0]), .in1(bm_d[7:0]), .in0(net295[0:7]),
     .sp12_v_b({sp12_v_b_bot[14], sp12_v_b_bot[12], sp12_v_b_bot[10],
     sp12_v_b_bot[8], sp12_v_b_bot[22], sp12_v_b_bot[6],
     sp12_v_b_bot[20], sp12_v_b_bot[4], sp12_v_b_bot[18],
     sp12_v_b_bot[2], sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_t ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}),
     .bl(bl[41:26]), .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12],
     sp12_v_b_top[10], sp12_v_b_top[8], sp12_v_b_top[22],
     sp12_v_b_top[6], sp12_v_b_top[20], sp12_v_b_top[4],
     sp12_v_b_top[18], sp12_v_b_top[2], sp12_v_b_top[16],
     sp12_v_b_top[0]}), .wl({wl_top[14], wl_top[15], wl_top[12],
     wl_top[13], wl_top[10], wl_top[11], wl_top[8], wl_top[9],
     wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2], wl_top[3],
     wl_top[0], wl_top[1]}), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .op(slf_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .sp12_h_r({sp12_h_r_top[22],
     sp12_h_r_top[6], sp12_h_r_top[20], sp12_h_r_top[4],
     sp12_h_r_top[18], sp12_h_r_top[2], sp12_h_r_top[16],
     sp12_h_r_top[0], sp12_h_r_top[14], sp12_h_r_top[12],
     sp12_h_r_top[10], sp12_h_r_top[8]}), .sp4_v_b({sp4_v_b_top[46],
     sp4_v_b_top[30], sp4_v_b_top[14], sp4_v_b_top[44],
     sp4_v_b_top[28], sp4_v_b_top[12], sp4_v_b_top[42],
     sp4_v_b_top[26], sp4_v_b_top[10], sp4_v_b_top[40],
     sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38], sp4_v_b_top[22],
     sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20], sp4_v_b_top[4],
     sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2], sp4_v_b_top[32],
     sp4_v_b_top[16], sp4_v_b_top[0]}), .sp4_r_v_b({sp4_r_v_b_top[47],
     sp4_r_v_b_top[31], sp4_r_v_b_top[15], sp4_r_v_b_top[45],
     sp4_r_v_b_top[29], sp4_r_v_b_top[13], sp4_r_v_b_top[43],
     sp4_r_v_b_top[27], sp4_r_v_b_top[11], sp4_r_v_b_top[41],
     sp4_r_v_b_top[25], sp4_r_v_b_top[9], sp4_r_v_b_top[39],
     sp4_r_v_b_top[23], sp4_r_v_b_top[7], sp4_r_v_b_top[37],
     sp4_r_v_b_top[21], sp4_r_v_b_top[5], sp4_r_v_b_top[35],
     sp4_r_v_b_top[19], sp4_r_v_b_top[3], sp4_r_v_b_top[33],
     sp4_r_v_b_top[17], sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46],
     sp4_h_r_top[30], sp4_h_r_top[14], sp4_h_r_top[44],
     sp4_h_r_top[28], sp4_h_r_top[12], sp4_h_r_top[42],
     sp4_h_r_top[26], sp4_h_r_top[10], sp4_h_r_top[40],
     sp4_h_r_top[24], sp4_h_r_top[8], sp4_h_r_top[38], sp4_h_r_top[22],
     sp4_h_r_top[6], sp4_h_r_top[36], sp4_h_r_top[20], sp4_h_r_top[4],
     sp4_h_r_top[34], sp4_h_r_top[18], sp4_h_r_top[2], sp4_h_r_top[32],
     sp4_h_r_top[16], sp4_h_r_top[0]}), .in3(bm_bweb[15:8]),
     .in2(in2_top[7:0]), .in1(bm_d[15:8]), .in0(net316[0:7]));

endmodule
// Library - leafcell, Cell - ice1f_array_BRAM_top, View - schematic
// LAST TIME SAVED: Feb 12 17:40:06 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module ice1f_array_BRAM_top ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, glb_netwk_bot, glb_netwk_top, slf_op_01,
     slf_op_02, slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07,
     slf_op_08, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02, sp4_h_l_03,
     sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07, sp4_h_l_08,
     sp4_h_r_01, sp4_h_r_02, sp4_h_r_03, sp4_h_r_04, sp4_h_r_05,
     sp4_h_r_06, sp4_h_r_07, sp4_h_r_08, sp4_r_v_b_01, sp4_r_v_b_02,
     sp4_r_v_b_03, sp4_r_v_b_04, sp4_r_v_b_05, sp4_r_v_b_06,
     sp4_r_v_b_07, sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03,
     sp4_v_b_04, sp4_v_b_05, sp4_v_b_06, sp4_v_b_07, sp4_v_b_08,
     sp4_v_t_08, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04,
     sp12_h_l_05, sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_r_01,
     sp12_h_r_02, sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06,
     sp12_h_r_07, sp12_h_r_08, sp12_v_b_01, sp12_v_t_08, vdd_cntl, wl,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i,
     bnl_op_01, bnr_op_01, bot_op_01, glb_netwk_col, lft_op_01,
     lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06, lft_op_07,
     lft_op_08, prog, rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04,
     rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, tnl_op_08, tnr_op_08,
     top_op_08 );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  slf_op_08;
output [7:0]  slf_op_04;
output [7:0]  slf_op_06;
output [7:0]  slf_op_02;
output [7:0]  slf_op_05;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_03;
output [7:0]  slf_op_07;
output [7:0]  slf_op_01;
output [7:0]  glb_netwk_bot;
output [7:0]  glb_netwk_top;

inout [47:0]  sp4_h_l_04;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_v_b_05;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_h_l_02;
inout [23:0]  sp12_h_l_04;
inout [47:0]  sp4_h_l_06;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_r_v_b_01;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_h_l_07;
inout [47:0]  sp4_r_v_b_04;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_h_r_01;
inout [23:0]  sp12_h_l_05;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_r_v_b_02;
inout [47:0]  sp4_h_l_03;
inout [23:0]  sp12_h_r_04;
inout [23:0]  sp12_v_t_08;
inout [47:0]  sp4_h_r_08;
inout [47:0]  sp4_v_b_07;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_h_r_05;
inout [23:0]  sp12_h_l_06;
inout [47:0]  sp4_h_r_04;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_r_v_b_05;
inout [47:0]  sp4_v_b_03;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_v_t_08;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_v_b_08;
inout [23:0]  sp12_h_r_03;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_r_v_b_03;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_h_l_08;
inout [47:0]  sp4_h_l_01;
inout [23:0]  sp12_h_r_08;
inout [47:0]  sp4_h_l_05;
inout [127:0]  reset_b;
inout [127:0]  wl;
inout [127:0]  vdd_cntl;
inout [23:0]  sp12_v_b_01;
inout [127:0]  pgate;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_v_b_06;

input [7:0]  rgt_op_01;
input [7:0]  tnl_op_08;
input [7:0]  bm_sa_i;
input [7:0]  rgt_op_02;
input [7:0]  lft_op_07;
input [7:0]  rgt_op_04;
input [7:0]  lft_op_02;
input [7:0]  lft_op_08;
input [7:0]  rgt_op_07;
input [7:0]  lft_op_03;
input [7:0]  rgt_op_06;
input [7:0]  bnr_op_01;
input [7:0]  glb_netwk_col;
input [7:0]  top_op_08;
input [7:0]  rgt_op_08;
input [7:0]  lft_op_05;
input [7:0]  bot_op_01;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_04;
input [7:0]  tnr_op_08;
input [7:0]  rgt_op_05;
input [7:0]  bnl_op_01;
input [7:0]  lft_op_01;
input [7:0]  lft_op_06;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net544;

wire  [0:7]  net481;

wire  [0:23]  net455;

wire  [7:0]  colbuf_cntl_top;

wire  [7:0]  colbuf_cntl_bot;

wire  [0:23]  net581;

wire  [0:23]  net518;

wire  [0:7]  net607;



clk_colbuf1kx8 I_clk_colbuf12kx8_b (
     .colbuf_cntl(colbuf_cntl_bot[7:0]), .col_clk(glb_netwk_bot[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_colbuf1kx8 I_clk_colbuf12kx8_t (
     .colbuf_cntl(colbuf_cntl_top[7:0]), .col_clk(glb_netwk_top[7:0]),
     .clk_in(glb_netwk_col[7:0]));
bram_4kprouting_tbankin I_bram_1516_in ( .bm_sdo_o(net491),
     .bm_sdi_i(net493), .bm_sclkrw_i(net494), .bm_sdo_i(bm_sdo_i),
     .bm_sweb_i(net495), .bm_sdi_o(bm_sdi_o),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_sweb_o(bm_sweb_o),
     .slf_op_top(slf_op_08[7:0]), .slf_op_bot(slf_op_07[7:0]),
     .wl_bot(wl[111:96]), .top_op_top(top_op_08[7:0]),
     .sp12_h_l_bot(sp12_h_l_07[23:0]), .sp4_h_l_bot(sp4_h_l_07[47:0]),
     .tnl_op_top(tnl_op_08[7:0]), .tnl_op_bot(lft_op_08[7:0]),
     .reset_b_top(reset_b[127:112]), .reset_b_bot(reset_b[111:96]),
     .vdd_cntl_top(vdd_cntl[127:112]), .prog(prog),
     .pgate_top(pgate[127:112]), .pgate_bot(pgate[111:96]),
     .lft_op_bot(lft_op_07[7:0]), .glb_netwk(glb_netwk_top[7:0]),
     .bm_wdummymux_en_i(net547), .bot_op_bot(slf_op_06[7:0]),
     .rgt_op_bot(rgt_op_07[7:0]), .bnl_op_top(lft_op_07[7:0]),
     .bnl_op_bot(lft_op_06[7:0]), .sp4_h_r_top(sp4_h_r_08[47:0]),
     .sp12_v_t_top(sp12_v_t_08[23:0]), .sp12_v_b_bot(net518[0:23]),
     .bm_init_i(net543), .sp4_h_r_bot(sp4_h_r_07[47:0]),
     .sp12_h_r_bot(sp12_h_r_07[23:0]), .sp4_v_t_top(sp4_v_t_08[47:0]),
     .sp4_v_b_bot(sp4_v_b_07[47:0]), .sp12_h_r_top(sp12_h_r_08[23:0]),
     .tnr_op_bot(rgt_op_08[7:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(net542), .sp4_h_l_top(sp4_h_l_08[47:0]),
     .lft_op_top(lft_op_08[7:0]), .wl_top(wl[127:112]),
     .sp12_h_l_top(sp12_h_l_08[23:0]), .sp4_v_b_top(sp4_v_b_08[47:0]),
     .tnr_op_top(tnr_op_08[7:0]), .rgt_op_top(rgt_op_08[7:0]),
     .bm_sa_i(net544[0:7]), .bm_sclk_i(net545), .bm_sreb_i(net546),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .vdd_cntl_bot(vdd_cntl[111:96]), .bnr_op_bot(rgt_op_06[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_07[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_08[47:0]), .bnr_op_top(rgt_op_07[7:0]));
bram_4kprouting_tbankout I_bram_out_0910 ( .bm_sdo_o(bm_sdo_o),
     .bm_sdi_i(bm_sdi_i), .bm_sclkrw_i(bm_sclkrw_i), .bm_sdo_i(net428),
     .bm_sweb_i(bm_sweb_i), .bm_sdi_o(net430), .bm_sclkrw_o(net431),
     .bm_sweb_o(net432), .slf_op_top(slf_op_02[7:0]),
     .slf_op_bot(slf_op_01[7:0]), .wl_top(wl[31:16]),
     .wl_bot(wl[15:0]), .top_op_top(slf_op_03[7:0]),
     .tnl_op_top(lft_op_03[7:0]), .tnl_op_bot(lft_op_02[7:0]),
     .reset_b_top(reset_b[31:16]), .reset_b_bot(reset_b[15:0]),
     .prog(prog), .pgate_top(pgate[31:16]), .pgate_bot(pgate[15:0]),
     .lft_op_top(lft_op_02[7:0]), .lft_op_bot(lft_op_01[7:0]),
     .glb_netwk(glb_netwk_bot[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bot_op_bot(bot_op_01[7:0]), .sp4_h_r_top(sp4_h_r_02[47:0]),
     .bnl_op_top(lft_op_01[7:0]), .bnl_op_bot(bnl_op_01[7:0]),
     .bnr_op_bot(bnr_op_01[7:0]), .sp4_h_r_bot(sp4_h_r_01[47:0]),
     .sp12_v_t_top(net455[0:23]), .sp12_v_b_bot(sp12_v_b_01[23:0]),
     .bm_init_i(bm_init_i), .sp12_h_l_top(sp12_h_l_02[23:0]),
     .sp12_h_r_bot(sp12_h_r_01[23:0]),
     .sp12_h_l_bot(sp12_h_l_01[23:0]),
     .sp12_h_r_top(sp12_h_r_02[23:0]), .sp4_v_t_top(sp4_v_b_03[47:0]),
     .sp4_v_b_top(sp4_v_b_02[47:0]), .sp4_v_b_bot(sp4_v_b_01[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_01[47:0]),
     .sp4_h_l_top(sp4_h_l_02[47:0]), .tnr_op_top(rgt_op_03[7:0]),
     .sp4_h_l_bot(sp4_h_l_01[47:0]), .tnr_op_bot(rgt_op_02[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .sp4_r_v_b_top(sp4_r_v_b_02[47:0]), .rgt_op_bot(rgt_op_01[7:0]),
     .rgt_op_top(rgt_op_02[7:0]), .bnr_op_top(rgt_op_01[7:0]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sreb_i(bm_sreb_i), .bm_rcapmux_en_o(net479),
     .bm_init_o(net480), .bm_sa_o(net481[0:7]), .bm_sclk_o(net482),
     .bm_sreb_o(net483), .bm_wdummymux_en_o(net484),
     .vdd_cntl_top(vdd_cntl[31:16]), .vdd_cntl_bot(vdd_cntl[15:0]));
bram_4kprouting_tbank I_bram_1314 (
     .cbit_colcntl(colbuf_cntl_top[7:0]), .bm_sdo_o(net554),
     .bm_sdi_i(net556), .bm_sclkrw_i(net557), .bm_sdo_i(net491),
     .bm_sweb_i(net558), .bm_sdi_o(net493), .bm_sclkrw_o(net494),
     .bm_sweb_o(net495), .slf_op_top(slf_op_06[7:0]),
     .slf_op_bot(slf_op_05[7:0]), .wl_top(wl[95:80]),
     .wl_bot(wl[79:64]), .top_op_top(slf_op_07[7:0]),
     .tnl_op_top(lft_op_07[7:0]), .tnl_op_bot(lft_op_06[7:0]),
     .reset_b_top(reset_b[95:80]), .reset_b_bot(reset_b[79:64]),
     .prog(prog), .pgate_top(pgate[95:80]), .pgate_bot(pgate[79:64]),
     .lft_op_top(lft_op_06[7:0]), .lft_op_bot(lft_op_05[7:0]),
     .glb_netwk(glb_netwk_top[7:0]), .bm_wdummymux_en_i(net610),
     .bot_op_bot(slf_op_04[7:0]), .sp4_h_r_top(sp4_h_r_06[47:0]),
     .bnl_op_top(lft_op_05[7:0]), .bnl_op_bot(lft_op_04[7:0]),
     .bnr_op_bot(rgt_op_04[7:0]), .sp4_h_r_bot(sp4_h_r_05[47:0]),
     .sp12_v_t_top(net518[0:23]), .sp12_v_b_bot(net581[0:23]),
     .bm_init_i(net606), .sp12_h_l_top(sp12_h_l_06[23:0]),
     .sp12_h_r_bot(sp12_h_r_05[23:0]),
     .sp12_h_l_bot(sp12_h_l_05[23:0]),
     .sp12_h_r_top(sp12_h_r_06[23:0]), .sp4_v_t_top(sp4_v_b_07[47:0]),
     .sp4_v_b_top(sp4_v_b_06[47:0]), .sp4_v_b_bot(sp4_v_b_05[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_05[47:0]),
     .sp4_h_l_top(sp4_h_l_06[47:0]), .tnr_op_top(rgt_op_07[7:0]),
     .sp4_h_l_bot(sp4_h_l_05[47:0]), .tnr_op_bot(rgt_op_06[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net605),
     .sp4_r_v_b_top(sp4_r_v_b_06[47:0]), .rgt_op_bot(rgt_op_05[7:0]),
     .rgt_op_top(rgt_op_06[7:0]), .bnr_op_top(rgt_op_05[7:0]),
     .bm_sa_i(net607[0:7]), .bm_sclk_i(net608), .bm_sreb_i(net609),
     .bm_rcapmux_en_o(net542), .bm_init_o(net543),
     .bm_sa_o(net544[0:7]), .bm_sclk_o(net545), .bm_sreb_o(net546),
     .bm_wdummymux_en_o(net547), .vdd_cntl_top(vdd_cntl[95:80]),
     .vdd_cntl_bot(vdd_cntl[79:64]));
bram_4kprouting_tbank I_bram_1112 (
     .cbit_colcntl(colbuf_cntl_bot[7:0]), .bm_sdo_o(net428),
     .bm_sdi_i(net430), .bm_sclkrw_i(net431), .bm_sdo_i(net554),
     .bm_sweb_i(net432), .bm_sdi_o(net556), .bm_sclkrw_o(net557),
     .bm_sweb_o(net558), .slf_op_top(slf_op_04[7:0]),
     .slf_op_bot(slf_op_03[7:0]), .wl_top(wl[63:48]),
     .wl_bot(wl[47:32]), .top_op_top(slf_op_05[7:0]),
     .tnl_op_top(lft_op_05[7:0]), .tnl_op_bot(lft_op_04[7:0]),
     .reset_b_top(reset_b[63:48]), .reset_b_bot(reset_b[47:32]),
     .prog(prog), .pgate_top(pgate[63:48]), .pgate_bot(pgate[47:32]),
     .lft_op_top(lft_op_04[7:0]), .lft_op_bot(lft_op_03[7:0]),
     .glb_netwk(glb_netwk_bot[7:0]), .bm_wdummymux_en_i(net484),
     .bot_op_bot(slf_op_02[7:0]), .sp4_h_r_top(sp4_h_r_04[47:0]),
     .bnl_op_top(lft_op_03[7:0]), .bnl_op_bot(lft_op_02[7:0]),
     .bnr_op_bot(rgt_op_02[7:0]), .sp4_h_r_bot(sp4_h_r_03[47:0]),
     .sp12_v_t_top(net581[0:23]), .sp12_v_b_bot(net455[0:23]),
     .bm_init_i(net480), .sp12_h_l_top(sp12_h_l_04[23:0]),
     .sp12_h_r_bot(sp12_h_r_03[23:0]),
     .sp12_h_l_bot(sp12_h_l_03[23:0]),
     .sp12_h_r_top(sp12_h_r_04[23:0]), .sp4_v_t_top(sp4_v_b_05[47:0]),
     .sp4_v_b_top(sp4_v_b_04[47:0]), .sp4_v_b_bot(sp4_v_b_03[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_03[47:0]),
     .sp4_h_l_top(sp4_h_l_04[47:0]), .tnr_op_top(rgt_op_05[7:0]),
     .sp4_h_l_bot(sp4_h_l_03[47:0]), .tnr_op_bot(rgt_op_04[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net479),
     .sp4_r_v_b_top(sp4_r_v_b_04[47:0]), .rgt_op_bot(rgt_op_03[7:0]),
     .rgt_op_top(rgt_op_04[7:0]), .bnr_op_top(rgt_op_03[7:0]),
     .bm_sa_i(net481[0:7]), .bm_sclk_i(net482), .bm_sreb_i(net483),
     .bm_rcapmux_en_o(net605), .bm_init_o(net606),
     .bm_sa_o(net607[0:7]), .bm_sclk_o(net608), .bm_sreb_o(net609),
     .bm_wdummymux_en_o(net610), .vdd_cntl_top(vdd_cntl[63:48]),
     .vdd_cntl_bot(vdd_cntl[47:32]));

endmodule
// Library - leafcell, Cell - ice1f_quad_tr, View - schematic
// LAST TIME SAVED: Jul 22 09:36:07 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module ice1f_quad_tr ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, ceb_o, cf_r, cf_t, fabric_out_07_17,
     fabric_out_08_17, fabric_out_13_09, fabric_out_13_10, hiz_b_o,
     mode_o, padeb_r, padeb_t_r, padin_07_17a, padin_13_09a, pado_r,
     pado_t_r, r_o, sdo, shift_o, slf_op_07_09, slf_op_07_10,
     slf_op_07_11, slf_op_07_12, slf_op_07_13, slf_op_07_14,
     slf_op_07_15, slf_op_07_16, slf_op_07_17, slf_op_08_09,
     slf_op_09_09, slf_op_10_09, slf_op_11_09, slf_op_12_09,
     slf_op_13_09, spi_ss_in_r_t, tclk_o, update_o, bl, pgate_r,
     reset_b_r, sp4_h_l_07_09, sp4_h_l_07_10, sp4_h_l_07_11,
     sp4_h_l_07_12, sp4_h_l_07_13, sp4_h_l_07_14, sp4_h_l_07_15,
     sp4_h_l_07_16, sp4_h_l_07_17, sp4_h_r_13_09, sp4_v_b_07_09,
     sp4_v_b_07_10, sp4_v_b_07_11, sp4_v_b_07_12, sp4_v_b_07_13,
     sp4_v_b_07_14, sp4_v_b_07_15, sp4_v_b_07_16, sp4_v_b_08_09,
     sp4_v_b_09_09, sp4_v_b_10_09, sp4_v_b_11_09, sp4_v_b_12_09,
     sp12_h_l_07_09, sp12_h_l_07_10, sp12_h_l_07_11, sp12_h_l_07_12,
     sp12_h_l_07_13, sp12_h_l_07_14, sp12_h_l_07_15, sp12_h_l_07_16,
     sp12_v_b_07_09, sp12_v_b_08_09, sp12_v_b_09_09, sp12_v_b_10_09,
     sp12_v_b_11_09, sp12_v_b_12_09, vdd_cntl_r, wl_r, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_07_09,
     bnl_op_08_09, bnl_op_09_09, bnl_op_10_09, bnl_op_11_09,
     bnl_op_12_09, bnl_op_13_09, bnr_op_07_09, bnr_op_08_09,
     bnr_op_09_09, bnr_op_10_09, bnr_op_11_09, bnr_op_12_09,
     bot_op_07_09, bot_op_08_09, bot_op_09_09, bot_op_10_09,
     bot_op_11_09, bot_op_12_09, bs_en_i, carry_in_07_09,
     carry_in_08_09, carry_in_09_09, carry_in_11_09, carry_in_12_09,
     ceb_i, end_of_startup_rgt_t, end_of_startup_top_r, glb_in,
     hiz_b_i, hold_r_t, hold_t_r, lft_op_07_09, lft_op_07_10,
     lft_op_07_11, lft_op_07_12, lft_op_07_13, lft_op_07_14,
     lft_op_07_15, lft_op_07_16, mode_i, padin_r, padin_t_r, prog,
     purst, r_i, sdi, shift_i, tclk_i, tiegnd, tievdd, tnl_op_07_16,
     update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bs_en_o, ceb_o,
     fabric_out_07_17, fabric_out_08_17, fabric_out_13_09,
     fabric_out_13_10, hiz_b_o, mode_o, padin_07_17a, padin_13_09a,
     r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en_i,
     carry_in_07_09, carry_in_08_09, carry_in_09_09, carry_in_11_09,
     carry_in_12_09, ceb_i, hiz_b_i, hold_r_t, hold_t_r, mode_i, prog,
     purst, r_i, sdi, shift_i, tclk_i, tiegnd, tievdd, update_i;

output [11:0]  padeb_r;
output [7:0]  slf_op_08_09;
output [7:0]  slf_op_07_16;
output [7:0]  slf_op_07_09;
output [7:0]  slf_op_11_09;
output [7:0]  slf_op_07_10;
output [7:0]  slf_op_07_11;
output [143:0]  cf_t;
output [7:0]  slf_op_07_14;
output [7:0]  slf_op_12_09;
output [11:0]  pado_t_r;
output [3:0]  slf_op_13_09;
output [7:0]  slf_op_09_09;
output [7:0]  slf_op_07_12;
output [15:0]  spi_ss_in_r_t;
output [7:0]  slf_op_07_13;
output [7:0]  slf_op_10_09;
output [191:0]  cf_r;
output [11:0]  padeb_t_r;
output [7:0]  slf_op_07_15;
output [3:0]  slf_op_07_17;
output [7:0]  bm_sa_o;
output [11:0]  pado_r;

inout [47:0]  sp4_h_l_07_14;
inout [23:0]  sp12_h_l_07_09;
inout [47:0]  sp4_v_b_07_11;
inout [23:0]  sp12_v_b_10_09;
inout [15:0]  sp4_h_r_13_09;
inout [23:0]  sp12_h_l_07_15;
inout [23:0]  sp12_h_l_07_14;
inout [23:0]  sp12_v_b_11_09;
inout [23:0]  sp12_v_b_09_09;
inout [47:0]  sp4_v_b_09_09;
inout [23:0]  sp12_h_l_07_12;
inout [47:0]  sp4_h_l_07_11;
inout [47:0]  sp4_v_b_10_09;
inout [47:0]  sp4_v_b_07_13;
inout [47:0]  sp4_v_b_07_10;
inout [23:0]  sp12_h_l_07_16;
inout [143:0]  vdd_cntl_r;
inout [47:0]  sp4_v_b_07_15;
inout [47:0]  sp4_v_b_07_12;
inout [47:0]  sp4_h_l_07_09;
inout [23:0]  sp12_h_l_07_10;
inout [47:0]  sp4_v_b_08_09;
inout [47:0]  sp4_v_b_07_09;
inout [23:0]  sp12_v_b_07_09;
inout [47:0]  sp4_h_l_07_12;
inout [23:0]  sp12_v_b_12_09;
inout [23:0]  sp12_v_b_08_09;
inout [47:0]  sp4_h_l_07_10;
inout [47:0]  sp4_v_b_11_09;
inout [15:0]  sp4_h_l_07_17;
inout [47:0]  sp4_v_b_07_14;
inout [47:0]  sp4_h_l_07_15;
inout [143:0]  pgate_r;
inout [47:0]  sp4_v_b_07_16;
inout [143:0]  wl_r;
inout [47:0]  sp4_h_l_07_13;
inout [329:0]  bl;
inout [23:0]  sp12_h_l_07_13;
inout [47:0]  sp4_v_b_12_09;
inout [23:0]  sp12_h_l_07_11;
inout [47:0]  sp4_h_l_07_16;
inout [143:0]  reset_b_r;

input [7:0]  lft_op_07_11;
input [7:0]  glb_in;
input [7:0]  bnr_op_08_09;
input [7:0]  bnl_op_13_09;
input [7:0]  bnl_op_11_09;
input [7:0]  bnl_op_07_09;
input [7:0]  bm_sa_i;
input [7:0]  bnr_op_09_09;
input [7:0]  bot_op_09_09;
input [7:0]  bnl_op_12_09;
input [7:0]  bnr_op_07_09;
input [11:0]  padin_r;
input [7:0]  bot_op_07_09;
input [7:0]  bot_op_08_09;
input [7:0]  bot_op_11_09;
input [11:0]  padin_t_r;
input [7:0]  lft_op_07_12;
input [7:0]  bnl_op_09_09;
input [7:0]  bnl_op_10_09;
input [16:9]  end_of_startup_rgt_t;
input [7:0]  lft_op_07_14;
input [7:0]  lft_op_07_16;
input [7:0]  bnr_op_10_09;
input [7:0]  lft_op_07_13;
input [7:0]  bot_op_12_09;
input [7:0]  bnr_op_11_09;
input [7:0]  bnr_op_12_09;
input [7:0]  lft_op_07_15;
input [7:0]  lft_op_07_09;
input [7:0]  bnl_op_08_09;
input [7:0]  bot_op_10_09;
input [7:0]  lft_op_07_10;
input [6:1]  end_of_startup_top_r;
input [3:0]  tnl_op_07_16;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:23]  net1318;

wire  [0:47]  net1398;

wire  [0:23]  net1248;

wire  [0:47]  net866;

wire  [0:23]  net895;

wire  [0:47]  net1427;

wire  [0:7]  net907;

wire  [0:23]  net968;

wire  [0:23]  net1340;

wire  [0:47]  net1187;

wire  [0:47]  net1093;

wire  [0:23]  net852;

wire  [0:47]  net889;

wire  [0:23]  net1247;

wire  [0:7]  net1381;

wire  [0:7]  net910;

wire  [0:47]  net1457;

wire  [0:47]  net1395;

wire  [0:47]  net974;

wire  [0:47]  net927;

wire  [0:47]  net1374;

wire  [0:7]  net1009;

wire  [0:47]  net1420;

wire  [0:47]  net1067;

wire  [0:47]  net1162;

wire  [0:47]  net1069;

wire  [0:23]  net970;

wire  [0:7]  net908;

wire  [0:47]  net1253;

wire  [0:7]  net1145;

wire  [0:23]  net1341;

wire  [0:0]  padinlat_r;

wire  [0:47]  net1188;

wire  [0:47]  net1116;

wire  [0:47]  net870;

wire  [0:47]  net975;

wire  [0:47]  net1212;

wire  [0:47]  net1160;

wire  [0:47]  net1397;

wire  [0:47]  net1396;

wire  [0:7]  net1196;

wire  [0:47]  net980;

wire  [0:47]  net1460;

wire  [0:23]  net1112;

wire  [0:47]  net1350;

wire  [0:47]  net1165;

wire  [0:7]  net959;

wire  [0:47]  net1023;

wire  [0:47]  net1074;

wire  [0:23]  net1299;

wire  [0:47]  net1002;

wire  [0:47]  net1303;

wire  [0:23]  net1154;

wire  [0:47]  net871;

wire  [0:47]  net979;

wire  [0:23]  net1063;

wire  [0:47]  net1210;

wire  [0:47]  net1167;

wire  [0:23]  net1205;

wire  [0:7]  net1135;

wire  [0:23]  net1020;

wire  [0:47]  net1095;

wire  [0:23]  net1297;

wire  [0:23]  net1156;

wire  [0:23]  net1204;

wire  [3:0]  slf_op_13_16;

wire  [0:47]  net1094;

wire  [0:7]  net1100;

wire  [0:23]  net834;

wire  [0:47]  net888;

wire  [0:7]  net1321;

wire  [0:7]  net904;

wire  [3:0]  slf_op_23_17;

wire  [0:23]  net1113;

wire  [0:7]  net1031;

wire  [0:47]  net1428;

wire  [0:47]  net1000;

wire  [0:23]  net1343;

wire  [0:47]  net1166;

wire  [0:7]  net951;

wire  [0:7]  net1103;

wire  [0:23]  net1392;

wire  [0:23]  net1155;

wire  [0:23]  net857;

wire  [0:47]  net1119;

wire  [0:47]  net1118;

wire  [0:47]  net1072;

wire  [0:47]  net1373;

wire  [0:7]  net1217;

wire  [0:7]  net1310;

wire  [0:47]  net921;

wire  [0:7]  net916;

wire  [0:23]  net1225;

wire  [0:23]  net1300;

wire  [0:47]  net1352;

wire  [0:47]  net891;

wire  [0:47]  net922;

wire  [0:47]  net1254;

wire  [0:7]  net949;

wire  [0:47]  net947;

wire  [0:23]  net1039;

wire  [0:47]  net1073;

wire  [0:47]  net1071;

wire  [0:47]  net1426;

wire  [3:0]  slf_op_13_15;

wire  [0:47]  net1348;

wire  [0:47]  net832;

wire  [0:47]  net999;

wire  [0:47]  net1459;

wire  [0:47]  net1260;

wire  [0:23]  net969;

wire  [0:47]  net920;

wire  [0:7]  net1044;

wire  [0:23]  net1298;

wire  [0:7]  net938;

wire  [0:23]  net1021;

wire  [0:47]  net1417;

wire  [0:23]  net1018;

wire  [3:0]  slf_op_12_17;

wire  [0:7]  net1423;

wire  [0:47]  net976;

wire  [0:23]  net893;

wire  [0:47]  net1446;

wire  [0:23]  net1390;

wire  [0:47]  net1092;

wire  [0:47]  net1025;

wire  [0:47]  net1371;

wire  [0:47]  net1319;

wire  [0:47]  net1346;

wire  [0:47]  net919;

wire  [0:7]  net1438;

wire  [0:47]  net1351;

wire  [0:47]  net1372;

wire  [0:47]  net1418;

wire  [0:23]  net1249;

wire  [0:7]  net1052;

wire  [0:23]  net1393;

wire  [3:0]  slf_op_40_17;

wire  [0:23]  net853;

wire  [3:0]  slf_op_13_12;

wire  [0:7]  net1422;

wire  [0:7]  net1431;

wire  [0:47]  net1164;

wire  [3:0]  slf_op_13_10;

wire  [0:7]  net1380;

wire  [0:23]  net1157;

wire  [0:23]  net946;

wire  [0:7]  net1430;

wire  [0:7]  net1195;

wire  [0:47]  net1117;

wire  [0:7]  net1137;

wire  [0:23]  net1342;

wire  [0:23]  net1114;

wire  [3:0]  slf_op_22_17;

wire  [0:7]  net1101;

wire  [0:23]  net1111;

wire  [0:7]  net1441;

wire  [0:23]  net1132;

wire  [0:7]  net1425;

wire  [0:23]  net1061;

wire  [0:47]  net1186;

wire  [0:23]  net1391;

wire  [0:47]  net1068;

wire  [0:7]  net1465;

wire  [3:0]  slf_op_13_14;

wire  [0:7]  net1042;

wire  [0:47]  net1353;

wire  [0:7]  net1435;

wire  [0:23]  net850;

wire  [3:0]  slf_op_13_13;

wire  [0:23]  net1207;

wire  [0:7]  net1010;

wire  [0:23]  net1250;

wire  [0:7]  net829;

wire  [0:47]  net1024;

wire  [0:47]  net1255;

wire  [0:47]  net1161;

wire  [0:7]  net917;

wire  [0:47]  net978;

wire  [0:47]  net1211;

wire  [0:23]  net1019;

wire  [0:47]  net1040;

wire  [0:23]  net854;

wire  [0:47]  net981;

wire  [0:47]  net873;

wire  [0:7]  net1323;

wire  [0:7]  net1124;

wire  [0:47]  net1026;

wire  [0:23]  net897;

wire  [0:47]  net868;

wire  [3:0]  slf_op_13_11;

wire  [0:7]  net1102;

wire  [0:47]  net890;

wire  [0:47]  net1421;

wire  [0:7]  net1008;

wire  [0:47]  net1133;

wire  [0:23]  net1206;

wire  [0:47]  net1001;

wire  [0:7]  net1424;

wire  [0:47]  net1185;

wire  [0:47]  net1347;

wire  [0:7]  net1331;

wire  [7:0]  clk_tree_drv;

wire  [0:23]  net1064;

wire  [0:23]  net1062;

wire  [0:7]  net1194;

wire  [0:15]  net776;

wire  [0:47]  net929;

wire  [0:23]  net971;

wire  [3:0]  slf_op_39_17;

wire  [0:0]  padinlat_t_r;

wire  [0:47]  net1209;

wire  [0:47]  net1226;

wire  [0:7]  net1382;



ice1f_array_RGT_IO_top12io I_preIO_rgt_t13 ( .padeb(padeb_r[11:0]),
     .pado(pado_r[11:0]), .padin(padin_r[11:0]),
     .cdone_in(end_of_startup_rgt_t[16:9]),
     .fabric_out_09(net_fabric_out_13_09),
     .fabric_out_10(net_fabric_out_13_10), .fabric_out_11(net691),
     .fabric_out_12(net692), .fabric_out_13(net693),
     .fabric_out_14(net694), .fabric_out_15(net695),
     .fabric_out_16(net696), .cf_r(cf_r[191:0]),
     .spi_ss_in_b(spi_ss_in_r_t[15:0]), .spiout({tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}), .spioeb({tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}),
     .wl(wl_r[127:0]), .vdd_cntl(vdd_cntl_r[127:0]),
     .reset_b(reset_b_r[127:0]), .pgate(pgate_r[127:0]),
     .SP4_h_l_13_16(net1428[0:47]), .SP12_h_l_13_16(net1300[0:23]),
     .lft_op_13_16(net1100[0:7]), .slf_op_13_16(slf_op_13_16[3:0]),
     .SP4_h_l_13_15(net1420[0:47]), .SP12_h_l_13_15(net1299[0:23]),
     .lft_op_13_15(net1101[0:7]), .slf_op_13_15(slf_op_13_15[3:0]),
     .SP4_h_l_13_14(net1427[0:47]), .SP12_h_l_13_14(net1298[0:23]),
     .lft_op_13_14(net1102[0:7]), .slf_op_13_14(slf_op_13_14[3:0]),
     .SP4_h_l_13_13(net1421[0:47]), .SP12_h_l_13_13(net1297[0:23]),
     .lft_op_13_13(net1103[0:7]), .slf_op_13_13(slf_op_13_13[3:0]),
     .SP4_h_l_13_12(net1426[0:47]), .SP12_h_l_13_12(net1247[0:23]),
     .lft_op_13_12(net1052[0:7]), .slf_op_13_12(slf_op_13_12[3:0]),
     .SP4_h_l_13_11(net1418[0:47]), .SP12_h_l_13_11(net1248[0:23]),
     .lft_op_13_11(net1042[0:7]), .slf_op_13_11(slf_op_13_11[3:0]),
     .SP4_h_l_13_10(net1417[0:47]), .SP12_h_l_13_10(net1249[0:23]),
     .lft_op_13_10(net1044[0:7]), .slf_op_13_10(slf_op_13_10[3:0]),
     .sp4_v_b_13_09(sp4_h_r_13_09[15:0]),
     .bnl_op_13_09(bnl_op_13_09[7:0]), .SP4_h_l_13_09(net1260[0:47]),
     .SP12_h_l_13_09(net1250[0:23]), .lft_op_13_09(slf_op_12_09[7:0]),
     .slf_op_13_09(slf_op_13_09[3:0]), .sp4_v_t_41_40(net776[0:15]),
     .tnl_op_41_40({slf_op_40_17[3], slf_op_40_17[2], slf_op_40_17[1],
     slf_op_40_17[0], slf_op_40_17[3], slf_op_40_17[2],
     slf_op_40_17[1], slf_op_40_17[0]}), .shift(shift_i),
     .bs_en(bs_en_i), .mode(mode_i), .sdi(sdi), .hiz_b(hiz_b_i),
     .prog(prog), .hold(hold_r_t), .update(update_i),
     .glb_netwk_col(clk_tree_drv[7:0]), .r(r_i), .sdo(net751),
     .bl(bl[329:312]), .tclk(tclk_i), .ceb(ceb_i));
pinlatbuf12p I_pinlatbuf12p ( .pad_in(padin_t_r[0]),
     .icegate(hold_t_r), .cbit(cf_t[15]), .cout(padinlat_t_r[0]),
     .prog(prog));
pinlatbuf12p I_pinlatbuf12p_r ( .pad_in(padin_r[0]),
     .icegate(hold_r_t), .cbit(cf_r[15]), .cout(padinlat_r[0]),
     .prog(prog));
scanbuf1f I_scanbuf_tr ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(net751), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_tr_1), .tclk_o(tclk_tr_1), .shift_o(shift_tr_1),
     .sdo(sdio_tr1), .r_o(r_tr_1), .mode_o(mode_tr_1),
     .hiz_b_o(hiz_b_tr_1), .ceb_o(ceb_tr_1), .bs_en_o(bs_en_tr_1));
ice1f_array_TOP_IO_rgt I_preio_top_r ( .pado_t_r(pado_t_r[11:0]),
     .padeb_t_r(padeb_t_r[11:0]), .padin_t_r(padin_t_r[11:0]),
     .fabric_out_08_17(net_fabric_out_08_17),
     .fabric_out_07_17(net_fabric_out_07_17),
     .bnl_op_07_17(lft_op_07_16[7:0]), .cf_top_l(cf_t[143:0]),
     .end_of_startup_top_l(end_of_startup_top_r[6:1]),
     .glb_net_11(net1031[0:7]), .glb_net_08(net938[0:7]),
     .glb_net_09(net1310[0:7]), .glb_net_12(net1217[0:7]),
     .glb_net_07(net1124[0:7]), .bl_07(bl[53:0]), .bl_08(bl[107:54]),
     .bl_09(bl[161:108]), .bl_11(bl[257:204]), .bl_12(bl[311:258]),
     .sp4_h_l_07_17(sp4_h_l_07_17[15:0]), .bl_10(bl[203:162]),
     .sp4_v_b_10_17(net832[0:47]), .sp4_h_r_12_17(net776[0:15]),
     .bnr_op_12_17({slf_op_13_16[3], slf_op_13_16[2], slf_op_13_16[1],
     slf_op_13_16[0], slf_op_13_16[3], slf_op_13_16[2],
     slf_op_13_16[1], slf_op_13_16[0]}), .sp4_v_b_07_17(net1133[0:47]),
     .slf_op_07_17(slf_op_07_17[3:0]),
     .lft_op_07_17(slf_op_07_16[7:0]), .sp12_v_b_07_17(net1132[0:23]),
     .sp4_v_b_08_17(net947[0:47]), .slf_op_08_17(slf_op_22_17[3:0]),
     .lft_op_08_17(net1430[0:7]), .sp12_v_b_08_17(net946[0:23]),
     .sp4_v_b_09_17(net1319[0:47]), .slf_op_09_17(slf_op_23_17[3:0]),
     .lft_op_09_17(net1438[0:7]), .sp12_v_b_09_17(net1318[0:23]),
     .slf_op_10_17(slf_op_12_17[3:0]), .lft_op_10_17(net1441[0:7]),
     .sp12_v_b_10_17(net834[0:23]), .sp4_v_b_11_17(net1040[0:47]),
     .slf_op_11_17(slf_op_39_17[3:0]), .lft_op_11_17(net1465[0:7]),
     .sp12_v_b_11_17(net1039[0:23]), .sp4_v_b_12_17(net1226[0:47]),
     .slf_op_12_17(slf_op_40_17[3:0]), .lft_op_12_17(net1100[0:7]),
     .sp12_v_b_12_17(net1225[0:23]), .hold_t_r(hold_t_r),
     .wl_l({wl_r[142], wl_r[143], wl_r[141], wl_r[140], wl_r[138],
     wl_r[139], wl_r[137], wl_r[136], wl_r[134], wl_r[135], wl_r[133],
     wl_r[132], wl_r[130], wl_r[131], wl_r[129], wl_r[128]}),
     .vdd_cntl_l({vdd_cntl_r[142], vdd_cntl_r[143], vdd_cntl_r[141],
     vdd_cntl_r[140], vdd_cntl_r[138], vdd_cntl_r[139],
     vdd_cntl_r[137], vdd_cntl_r[136], vdd_cntl_r[134],
     vdd_cntl_r[135], vdd_cntl_r[133], vdd_cntl_r[132],
     vdd_cntl_r[130], vdd_cntl_r[131], vdd_cntl_r[129],
     vdd_cntl_r[128]}), .update_i(update_tr_1), .tievdd(tievdd),
     .tiegnd(tiegnd), .tclk_i(tclk_tr_1), .shift_i(shift_tr_1),
     .sdi(sdio_tr1), .reset_l({reset_b_r[142], reset_b_r[143],
     reset_b_r[141], reset_b_r[140], reset_b_r[138], reset_b_r[139],
     reset_b_r[137], reset_b_r[136], reset_b_r[134], reset_b_r[135],
     reset_b_r[133], reset_b_r[132], reset_b_r[130], reset_b_r[131],
     reset_b_r[129], reset_b_r[128]}), .r_i(r_tr_1), .prog(prog),
     .pgate_l({pgate_r[142], pgate_r[143], pgate_r[141], pgate_r[140],
     pgate_r[138], pgate_r[139], pgate_r[137], pgate_r[136],
     pgate_r[134], pgate_r[135], pgate_r[133], pgate_r[132],
     pgate_r[130], pgate_r[131], pgate_r[129], pgate_r[128]}),
     .mode_i(mode_tr_1), .hiz_b_i(hiz_b_tr_1), .bs_en_i(bs_en_tr_1),
     .update_o(update_o), .tclk_o(tclk_o), .shift_o(shift_o),
     .sdo(sdo), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .glb_net_10(net829[0:7]), .bs_en_o(bs_en_o), .ceb_o(ceb_o),
     .ceb_i(ceb_tr_1));
ice1f_array_BRAM_top I_array_BRAM_t10 ( .glb_netwk_bot(net1422[0:7]),
     .glb_netwk_top(net829[0:7]), .tnr_op_08({slf_op_39_17[3],
     slf_op_39_17[2], slf_op_39_17[1], slf_op_39_17[0],
     slf_op_39_17[3], slf_op_39_17[2], slf_op_39_17[1],
     slf_op_39_17[0]}), .tnl_op_08({slf_op_23_17[3], slf_op_23_17[2],
     slf_op_23_17[1], slf_op_23_17[0], slf_op_23_17[3],
     slf_op_23_17[2], slf_op_23_17[1], slf_op_23_17[0]}),
     .sp4_v_t_08(net832[0:47]), .top_op_08({slf_op_12_17[3],
     slf_op_12_17[2], slf_op_12_17[1], slf_op_12_17[0],
     slf_op_12_17[3], slf_op_12_17[2], slf_op_12_17[1],
     slf_op_12_17[0]}), .sp12_v_t_08(net834[0:23]),
     .pgate(pgate_r[127:0]), .vdd_cntl(vdd_cntl_r[127:0]),
     .reset_b(reset_b_r[127:0]), .wl(wl_r[127:0]), .prog(prog),
     .glb_netwk_col(clk_tree_drv[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .sp12_h_l_07(net1392[0:23]), .sp4_v_b_08(net1398[0:47]),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bnr_op_01(bnr_op_10_09[7:0]), .sp12_h_r_06(net850[0:23]),
     .sp12_h_l_06(net1391[0:23]), .sp12_h_r_05(net852[0:23]),
     .sp12_h_r_08(net853[0:23]), .sp12_h_r_03(net854[0:23]),
     .sp12_h_l_08(net1393[0:23]), .sp12_h_l_05(net1390[0:23]),
     .sp12_h_r_07(net857[0:23]), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_sreb_o(bm_sreb_o), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .sp4_r_v_b_01(sp4_v_b_11_09[47:0]),
     .sp4_v_b_02(net1348[0:47]), .sp4_r_v_b_02(net866[0:47]),
     .sp4_v_b_03(net1347[0:47]), .sp4_r_v_b_03(net868[0:47]),
     .sp4_v_b_04(net1346[0:47]), .sp4_r_v_b_04(net870[0:47]),
     .sp4_r_v_b_06(net871[0:47]), .sp4_v_b_06(net1396[0:47]),
     .sp4_r_v_b_05(net873[0:47]), .sp4_v_b_05(net1395[0:47]),
     .lft_op_08(net1438[0:7]), .lft_op_07(net1008[0:7]),
     .lft_op_06(net1009[0:7]), .lft_op_05(net1010[0:7]),
     .sp4_v_b_07(net1397[0:47]), .sp12_h_l_03(net1341[0:23]),
     .sp12_h_l_04(net1340[0:23]), .sp12_h_l_02(net1342[0:23]),
     .sp12_h_l_01(net1343[0:23]), .slf_op_07(net1380[0:7]),
     .slf_op_08(net1441[0:7]), .sp4_h_l_07(net1372[0:47]),
     .sp4_h_l_08(net1371[0:47]), .sp4_h_r_07(net888[0:47]),
     .sp4_h_r_08(net889[0:47]), .sp4_r_v_b_07(net890[0:47]),
     .sp4_r_v_b_08(net891[0:47]), .sp4_v_b_01(sp4_v_b_10_09[47:0]),
     .sp12_h_r_01(net893[0:23]), .bm_sdo_i(bm_sdo_i),
     .sp12_h_r_02(net895[0:23]), .bl(bl[203:162]),
     .sp12_h_r_04(net897[0:23]), .sp12_v_b_01(sp12_v_b_10_09[23:0]),
     .bnl_op_01(bnl_op_10_09[7:0]), .lft_op_01(slf_op_09_09[7:0]),
     .lft_op_02(net951[0:7]), .lft_op_03(net949[0:7]),
     .lft_op_04(net959[0:7]), .rgt_op_07(net904[0:7]),
     .rgt_op_08(net1465[0:7]), .bot_op_01(bot_op_10_09[7:0]),
     .rgt_op_03(net907[0:7]), .rgt_op_02(net908[0:7]),
     .rgt_op_01(slf_op_11_09[7:0]), .rgt_op_04(net910[0:7]),
     .slf_op_04(net1331[0:7]), .slf_op_03(net1321[0:7]),
     .slf_op_02(net1323[0:7]), .slf_op_01(slf_op_10_09[7:0]),
     .slf_op_06(net1381[0:7]), .rgt_op_05(net916[0:7]),
     .rgt_op_06(net917[0:7]), .slf_op_05(net1382[0:7]),
     .sp4_h_r_04(net919[0:47]), .sp4_h_r_03(net920[0:47]),
     .sp4_h_r_02(net921[0:47]), .sp4_h_r_01(net922[0:47]),
     .sp4_h_l_04(net1350[0:47]), .sp4_h_l_03(net1351[0:47]),
     .sp4_h_l_02(net1352[0:47]), .sp4_h_l_01(net1353[0:47]),
     .sp4_h_r_06(net927[0:47]), .sp4_h_l_06(net1373[0:47]),
     .sp4_h_r_05(net929[0:47]), .sp4_h_l_05(net1374[0:47]),
     .bm_sdo_o(bm_sdo_o), .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_sweb_i(bm_sweb_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sweb_o(bm_sweb_o));
ice1f_array_LT_top I_lt_col_t08 ( .glb_netwk_to(net938[0:7]),
     .glb_netwk_bo(net1425[0:7]), .vdd_cntl(vdd_cntl_r[127:0]),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .top_op_08({slf_op_22_17[3], slf_op_22_17[2], slf_op_22_17[1],
     slf_op_22_17[0], slf_op_22_17[3], slf_op_22_17[2],
     slf_op_22_17[1], slf_op_22_17[0]}), .tnl_op_08({slf_op_07_17[3],
     slf_op_07_17[2], slf_op_07_17[1], slf_op_07_17[0],
     slf_op_07_17[3], slf_op_07_17[2], slf_op_07_17[1],
     slf_op_07_17[0]}), .tnr_op_08({slf_op_23_17[3], slf_op_23_17[2],
     slf_op_23_17[1], slf_op_23_17[0], slf_op_23_17[3],
     slf_op_23_17[2], slf_op_23_17[1], slf_op_23_17[0]}),
     .sp12_v_t_08(net946[0:23]), .sp4_v_t_08(net947[0:47]),
     .wl(wl_r[127:0]), .rgt_op_03(net949[0:7]),
     .slf_op_02(net1137[0:7]), .rgt_op_02(net951[0:7]),
     .rgt_op_01(slf_op_09_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(slf_op_07_12[7:0]), .lft_op_03(slf_op_07_11[7:0]),
     .lft_op_02(slf_op_07_10[7:0]), .lft_op_01(slf_op_07_09[7:0]),
     .rgt_op_04(net959[0:7]), .carry_in(carry_in_08_09),
     .bnl_op_01(bnl_op_08_09[7:0]), .slf_op_04(net1145[0:7]),
     .slf_op_03(net1135[0:7]), .slf_op_01(slf_op_08_09[7:0]),
     .sp4_h_l_04(net1164[0:47]), .carry_out(net966),
     .sp12_v_b__01(sp12_v_b_08_09[23:0]), .sp12_h_r_04(net968[0:23]),
     .sp12_h_r_03(net969[0:23]), .sp12_h_r_02(net970[0:23]),
     .sp12_h_r_01(net971[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_08_09[47:0]), .sp4_r_v_b_04(net974[0:47]),
     .sp4_r_v_b_03(net975[0:47]), .sp4_r_v_b_02(net976[0:47]),
     .sp4_r_v_b_01(sp4_v_b_09_09[47:0]), .sp4_h_r_04(net978[0:47]),
     .sp4_h_r_03(net979[0:47]), .sp4_h_r_02(net980[0:47]),
     .sp4_h_r_01(net981[0:47]), .sp4_h_l_03(net1165[0:47]),
     .sp4_h_l_02(net1166[0:47]), .sp4_h_l_01(net1167[0:47]),
     .bl(bl[107:54]), .bot_op_01(bot_op_08_09[7:0]),
     .sp12_h_l_01(net1157[0:23]), .sp12_h_l_02(net1156[0:23]),
     .sp12_h_l_03(net1155[0:23]), .sp12_h_l_04(net1154[0:23]),
     .sp4_v_b_04(net1160[0:47]), .sp4_v_b_03(net1161[0:47]),
     .sp4_v_b_02(net1162[0:47]), .bnr_op_01(bnr_op_08_09[7:0]),
     .sp4_h_l_05(net1188[0:47]), .sp4_h_l_06(net1187[0:47]),
     .sp4_h_l_07(net1186[0:47]), .sp4_h_l_08(net1185[0:47]),
     .sp4_h_r_08(net999[0:47]), .sp4_h_r_07(net1000[0:47]),
     .sp4_h_r_06(net1001[0:47]), .sp4_h_r_05(net1002[0:47]),
     .slf_op_05(net1196[0:7]), .slf_op_06(net1195[0:7]),
     .slf_op_07(net1194[0:7]), .slf_op_08(net1430[0:7]),
     .rgt_op_08(net1438[0:7]), .rgt_op_07(net1008[0:7]),
     .rgt_op_06(net1009[0:7]), .rgt_op_05(net1010[0:7]),
     .lft_op_08(slf_op_07_16[7:0]), .lft_op_07(slf_op_07_15[7:0]),
     .lft_op_06(slf_op_07_14[7:0]), .lft_op_05(slf_op_07_13[7:0]),
     .sp12_h_l_08(net1207[0:23]), .sp12_h_l_07(net1206[0:23]),
     .sp12_h_l_06(net1205[0:23]), .sp12_h_r_05(net1018[0:23]),
     .sp12_h_r_06(net1019[0:23]), .sp12_h_r_07(net1020[0:23]),
     .sp12_h_r_08(net1021[0:23]), .sp12_h_l_05(net1204[0:23]),
     .sp4_r_v_b_05(net1023[0:47]), .sp4_r_v_b_06(net1024[0:47]),
     .sp4_r_v_b_07(net1025[0:47]), .sp4_r_v_b_08(net1026[0:47]),
     .sp4_v_b_08(net1212[0:47]), .sp4_v_b_07(net1211[0:47]),
     .sp4_v_b_06(net1210[0:47]), .sp4_v_b_05(net1209[0:47]));
ice1f_array_LT_top I_lt_col_t11 ( .glb_netwk_to(net1031[0:7]),
     .glb_netwk_bo(net1431[0:7]), .vdd_cntl(vdd_cntl_r[127:0]),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .top_op_08({slf_op_39_17[3], slf_op_39_17[2], slf_op_39_17[1],
     slf_op_39_17[0], slf_op_39_17[3], slf_op_39_17[2],
     slf_op_39_17[1], slf_op_39_17[0]}), .tnl_op_08({slf_op_12_17[3],
     slf_op_12_17[2], slf_op_12_17[1], slf_op_12_17[0],
     slf_op_12_17[3], slf_op_12_17[2], slf_op_12_17[1],
     slf_op_12_17[0]}), .tnr_op_08({slf_op_40_17[3], slf_op_40_17[2],
     slf_op_40_17[1], slf_op_40_17[0], slf_op_40_17[3],
     slf_op_40_17[2], slf_op_40_17[1], slf_op_40_17[0]}),
     .sp12_v_t_08(net1039[0:23]), .sp4_v_t_08(net1040[0:47]),
     .wl(wl_r[127:0]), .rgt_op_03(net1042[0:7]),
     .slf_op_02(net908[0:7]), .rgt_op_02(net1044[0:7]),
     .rgt_op_01(slf_op_12_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net1331[0:7]), .lft_op_03(net1321[0:7]),
     .lft_op_02(net1323[0:7]), .lft_op_01(slf_op_10_09[7:0]),
     .rgt_op_04(net1052[0:7]), .carry_in(carry_in_11_09),
     .bnl_op_01(bnl_op_11_09[7:0]), .slf_op_04(net910[0:7]),
     .slf_op_03(net907[0:7]), .slf_op_01(slf_op_11_09[7:0]),
     .sp4_h_l_04(net919[0:47]), .carry_out(net1059),
     .sp12_v_b__01(sp12_v_b_11_09[23:0]), .sp12_h_r_04(net1061[0:23]),
     .sp12_h_r_03(net1062[0:23]), .sp12_h_r_02(net1063[0:23]),
     .sp12_h_r_01(net1064[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_11_09[47:0]), .sp4_r_v_b_04(net1067[0:47]),
     .sp4_r_v_b_03(net1068[0:47]), .sp4_r_v_b_02(net1069[0:47]),
     .sp4_r_v_b_01(sp4_v_b_12_09[47:0]), .sp4_h_r_04(net1071[0:47]),
     .sp4_h_r_03(net1072[0:47]), .sp4_h_r_02(net1073[0:47]),
     .sp4_h_r_01(net1074[0:47]), .sp4_h_l_03(net920[0:47]),
     .sp4_h_l_02(net921[0:47]), .sp4_h_l_01(net922[0:47]),
     .bl(bl[257:204]), .bot_op_01(bot_op_11_09[7:0]),
     .sp12_h_l_01(net893[0:23]), .sp12_h_l_02(net895[0:23]),
     .sp12_h_l_03(net854[0:23]), .sp12_h_l_04(net897[0:23]),
     .sp4_v_b_04(net870[0:47]), .sp4_v_b_03(net868[0:47]),
     .sp4_v_b_02(net866[0:47]), .bnr_op_01(bnr_op_11_09[7:0]),
     .sp4_h_l_05(net929[0:47]), .sp4_h_l_06(net927[0:47]),
     .sp4_h_l_07(net888[0:47]), .sp4_h_l_08(net889[0:47]),
     .sp4_h_r_08(net1092[0:47]), .sp4_h_r_07(net1093[0:47]),
     .sp4_h_r_06(net1094[0:47]), .sp4_h_r_05(net1095[0:47]),
     .slf_op_05(net916[0:7]), .slf_op_06(net917[0:7]),
     .slf_op_07(net904[0:7]), .slf_op_08(net1465[0:7]),
     .rgt_op_08(net1100[0:7]), .rgt_op_07(net1101[0:7]),
     .rgt_op_06(net1102[0:7]), .rgt_op_05(net1103[0:7]),
     .lft_op_08(net1441[0:7]), .lft_op_07(net1380[0:7]),
     .lft_op_06(net1381[0:7]), .lft_op_05(net1382[0:7]),
     .sp12_h_l_08(net853[0:23]), .sp12_h_l_07(net857[0:23]),
     .sp12_h_l_06(net850[0:23]), .sp12_h_r_05(net1111[0:23]),
     .sp12_h_r_06(net1112[0:23]), .sp12_h_r_07(net1113[0:23]),
     .sp12_h_r_08(net1114[0:23]), .sp12_h_l_05(net852[0:23]),
     .sp4_r_v_b_05(net1116[0:47]), .sp4_r_v_b_06(net1117[0:47]),
     .sp4_r_v_b_07(net1118[0:47]), .sp4_r_v_b_08(net1119[0:47]),
     .sp4_v_b_08(net891[0:47]), .sp4_v_b_07(net890[0:47]),
     .sp4_v_b_06(net871[0:47]), .sp4_v_b_05(net873[0:47]));
ice1f_array_LT_top I_lt_col_t07 ( .glb_netwk_to(net1124[0:7]),
     .glb_netwk_bo(net1423[0:7]), .vdd_cntl(vdd_cntl_r[127:0]),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .top_op_08({slf_op_07_17[3], slf_op_07_17[2], slf_op_07_17[1],
     slf_op_07_17[0], slf_op_07_17[3], slf_op_07_17[2],
     slf_op_07_17[1], slf_op_07_17[0]}), .tnl_op_08({tnl_op_07_16[3],
     tnl_op_07_16[2], tnl_op_07_16[1], tnl_op_07_16[0],
     tnl_op_07_16[3], tnl_op_07_16[2], tnl_op_07_16[1],
     tnl_op_07_16[0]}), .tnr_op_08({slf_op_22_17[3], slf_op_22_17[2],
     slf_op_22_17[1], slf_op_22_17[0], slf_op_22_17[3],
     slf_op_22_17[2], slf_op_22_17[1], slf_op_22_17[0]}),
     .sp12_v_t_08(net1132[0:23]), .sp4_v_t_08(net1133[0:47]),
     .wl(wl_r[127:0]), .rgt_op_03(net1135[0:7]),
     .slf_op_02(slf_op_07_10[7:0]), .rgt_op_02(net1137[0:7]),
     .rgt_op_01(slf_op_08_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(lft_op_07_12[7:0]), .lft_op_03(lft_op_07_11[7:0]),
     .lft_op_02(lft_op_07_10[7:0]), .lft_op_01(lft_op_07_09[7:0]),
     .rgt_op_04(net1145[0:7]), .carry_in(carry_in_07_09),
     .bnl_op_01(bnl_op_07_09[7:0]), .slf_op_04(slf_op_07_12[7:0]),
     .slf_op_03(slf_op_07_11[7:0]), .slf_op_01(slf_op_07_09[7:0]),
     .sp4_h_l_04(sp4_h_l_07_12[47:0]), .carry_out(net1432),
     .sp12_v_b__01(sp12_v_b_07_09[23:0]), .sp12_h_r_04(net1154[0:23]),
     .sp12_h_r_03(net1155[0:23]), .sp12_h_r_02(net1156[0:23]),
     .sp12_h_r_01(net1157[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_07_09[47:0]), .sp4_r_v_b_04(net1160[0:47]),
     .sp4_r_v_b_03(net1161[0:47]), .sp4_r_v_b_02(net1162[0:47]),
     .sp4_r_v_b_01(sp4_v_b_08_09[47:0]), .sp4_h_r_04(net1164[0:47]),
     .sp4_h_r_03(net1165[0:47]), .sp4_h_r_02(net1166[0:47]),
     .sp4_h_r_01(net1167[0:47]), .sp4_h_l_03(sp4_h_l_07_11[47:0]),
     .sp4_h_l_02(sp4_h_l_07_10[47:0]),
     .sp4_h_l_01(sp4_h_l_07_09[47:0]), .bl(bl[53:0]),
     .bot_op_01(bot_op_07_09[7:0]), .sp12_h_l_01(sp12_h_l_07_09[23:0]),
     .sp12_h_l_02(sp12_h_l_07_10[23:0]),
     .sp12_h_l_03(sp12_h_l_07_11[23:0]),
     .sp12_h_l_04(sp12_h_l_07_12[23:0]),
     .sp4_v_b_04(sp4_v_b_07_12[47:0]),
     .sp4_v_b_03(sp4_v_b_07_11[47:0]),
     .sp4_v_b_02(sp4_v_b_07_10[47:0]), .bnr_op_01(bnr_op_07_09[7:0]),
     .sp4_h_l_05(sp4_h_l_07_13[47:0]),
     .sp4_h_l_06(sp4_h_l_07_14[47:0]),
     .sp4_h_l_07(sp4_h_l_07_15[47:0]),
     .sp4_h_l_08(sp4_h_l_07_16[47:0]), .sp4_h_r_08(net1185[0:47]),
     .sp4_h_r_07(net1186[0:47]), .sp4_h_r_06(net1187[0:47]),
     .sp4_h_r_05(net1188[0:47]), .slf_op_05(slf_op_07_13[7:0]),
     .slf_op_06(slf_op_07_14[7:0]), .slf_op_07(slf_op_07_15[7:0]),
     .slf_op_08(slf_op_07_16[7:0]), .rgt_op_08(net1430[0:7]),
     .rgt_op_07(net1194[0:7]), .rgt_op_06(net1195[0:7]),
     .rgt_op_05(net1196[0:7]), .lft_op_08(lft_op_07_16[7:0]),
     .lft_op_07(lft_op_07_15[7:0]), .lft_op_06(lft_op_07_14[7:0]),
     .lft_op_05(lft_op_07_13[7:0]), .sp12_h_l_08(sp12_h_l_07_16[23:0]),
     .sp12_h_l_07(sp12_h_l_07_15[23:0]),
     .sp12_h_l_06(sp12_h_l_07_14[23:0]), .sp12_h_r_05(net1204[0:23]),
     .sp12_h_r_06(net1205[0:23]), .sp12_h_r_07(net1206[0:23]),
     .sp12_h_r_08(net1207[0:23]), .sp12_h_l_05(sp12_h_l_07_13[23:0]),
     .sp4_r_v_b_05(net1209[0:47]), .sp4_r_v_b_06(net1210[0:47]),
     .sp4_r_v_b_07(net1211[0:47]), .sp4_r_v_b_08(net1212[0:47]),
     .sp4_v_b_08(sp4_v_b_07_16[47:0]),
     .sp4_v_b_07(sp4_v_b_07_15[47:0]),
     .sp4_v_b_06(sp4_v_b_07_14[47:0]),
     .sp4_v_b_05(sp4_v_b_07_13[47:0]));
ice1f_array_LT_top I_lt_col_t12 ( .glb_netwk_to(net1217[0:7]),
     .glb_netwk_bo(net1435[0:7]), .vdd_cntl(vdd_cntl_r[127:0]),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .top_op_08({slf_op_40_17[3], slf_op_40_17[2], slf_op_40_17[1],
     slf_op_40_17[0], slf_op_40_17[3], slf_op_40_17[2],
     slf_op_40_17[1], slf_op_40_17[0]}), .tnl_op_08({slf_op_39_17[3],
     slf_op_39_17[2], slf_op_39_17[1], slf_op_39_17[0],
     slf_op_39_17[3], slf_op_39_17[2], slf_op_39_17[1],
     slf_op_39_17[0]}), .tnr_op_08({tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd}), .sp12_v_t_08(net1225[0:23]),
     .sp4_v_t_08(net1226[0:47]), .wl(wl_r[127:0]),
     .rgt_op_03({slf_op_13_11[3], slf_op_13_11[2], slf_op_13_11[1],
     slf_op_13_11[0], slf_op_13_11[3], slf_op_13_11[2],
     slf_op_13_11[1], slf_op_13_11[0]}), .slf_op_02(net1044[0:7]),
     .rgt_op_02({slf_op_13_10[3], slf_op_13_10[2], slf_op_13_10[1],
     slf_op_13_10[0], slf_op_13_10[3], slf_op_13_10[2],
     slf_op_13_10[1], slf_op_13_10[0]}), .rgt_op_01({slf_op_13_09[3],
     slf_op_13_09[2], slf_op_13_09[1], slf_op_13_09[0],
     slf_op_13_09[3], slf_op_13_09[2], slf_op_13_09[1],
     slf_op_13_09[0]}), .purst(purst), .prog(prog),
     .lft_op_04(net910[0:7]), .lft_op_03(net907[0:7]),
     .lft_op_02(net908[0:7]), .lft_op_01(slf_op_11_09[7:0]),
     .rgt_op_04({slf_op_13_12[3], slf_op_13_12[2], slf_op_13_12[1],
     slf_op_13_12[0], slf_op_13_12[3], slf_op_13_12[2],
     slf_op_13_12[1], slf_op_13_12[0]}), .carry_in(carry_in_12_09),
     .bnl_op_01(bnl_op_12_09[7:0]), .slf_op_04(net1052[0:7]),
     .slf_op_03(net1042[0:7]), .slf_op_01(slf_op_12_09[7:0]),
     .sp4_h_l_04(net1071[0:47]), .carry_out(net1245),
     .sp12_v_b__01(sp12_v_b_12_09[23:0]), .sp12_h_r_04(net1247[0:23]),
     .sp12_h_r_03(net1248[0:23]), .sp12_h_r_02(net1249[0:23]),
     .sp12_h_r_01(net1250[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_12_09[47:0]), .sp4_r_v_b_04(net1253[0:47]),
     .sp4_r_v_b_03(net1254[0:47]), .sp4_r_v_b_02(net1255[0:47]),
     .sp4_r_v_b_01(net1446[0:47]), .sp4_h_r_04(net1426[0:47]),
     .sp4_h_r_03(net1418[0:47]), .sp4_h_r_02(net1417[0:47]),
     .sp4_h_r_01(net1260[0:47]), .sp4_h_l_03(net1072[0:47]),
     .sp4_h_l_02(net1073[0:47]), .sp4_h_l_01(net1074[0:47]),
     .bl(bl[311:258]), .bot_op_01(bot_op_12_09[7:0]),
     .sp12_h_l_01(net1064[0:23]), .sp12_h_l_02(net1063[0:23]),
     .sp12_h_l_03(net1062[0:23]), .sp12_h_l_04(net1061[0:23]),
     .sp4_v_b_04(net1067[0:47]), .sp4_v_b_03(net1068[0:47]),
     .sp4_v_b_02(net1069[0:47]), .bnr_op_01(bnr_op_12_09[7:0]),
     .sp4_h_l_05(net1095[0:47]), .sp4_h_l_06(net1094[0:47]),
     .sp4_h_l_07(net1093[0:47]), .sp4_h_l_08(net1092[0:47]),
     .sp4_h_r_08(net1428[0:47]), .sp4_h_r_07(net1420[0:47]),
     .sp4_h_r_06(net1427[0:47]), .sp4_h_r_05(net1421[0:47]),
     .slf_op_05(net1103[0:7]), .slf_op_06(net1102[0:7]),
     .slf_op_07(net1101[0:7]), .slf_op_08(net1100[0:7]),
     .rgt_op_08({slf_op_13_16[3], slf_op_13_16[2], slf_op_13_16[1],
     slf_op_13_16[0], slf_op_13_16[3], slf_op_13_16[2],
     slf_op_13_16[1], slf_op_13_16[0]}), .rgt_op_07({slf_op_13_15[3],
     slf_op_13_15[2], slf_op_13_15[1], slf_op_13_15[0],
     slf_op_13_15[3], slf_op_13_15[2], slf_op_13_15[1],
     slf_op_13_15[0]}), .rgt_op_06({slf_op_13_14[3], slf_op_13_14[2],
     slf_op_13_14[1], slf_op_13_14[0], slf_op_13_14[3],
     slf_op_13_14[2], slf_op_13_14[1], slf_op_13_14[0]}),
     .rgt_op_05({slf_op_13_13[3], slf_op_13_13[2], slf_op_13_13[1],
     slf_op_13_13[0], slf_op_13_13[3], slf_op_13_13[2],
     slf_op_13_13[1], slf_op_13_13[0]}), .lft_op_08(net1465[0:7]),
     .lft_op_07(net904[0:7]), .lft_op_06(net917[0:7]),
     .lft_op_05(net916[0:7]), .sp12_h_l_08(net1114[0:23]),
     .sp12_h_l_07(net1113[0:23]), .sp12_h_l_06(net1112[0:23]),
     .sp12_h_r_05(net1297[0:23]), .sp12_h_r_06(net1298[0:23]),
     .sp12_h_r_07(net1299[0:23]), .sp12_h_r_08(net1300[0:23]),
     .sp12_h_l_05(net1111[0:23]), .sp4_r_v_b_05(net1459[0:47]),
     .sp4_r_v_b_06(net1303[0:47]), .sp4_r_v_b_07(net1457[0:47]),
     .sp4_r_v_b_08(net1460[0:47]), .sp4_v_b_08(net1119[0:47]),
     .sp4_v_b_07(net1118[0:47]), .sp4_v_b_06(net1117[0:47]),
     .sp4_v_b_05(net1116[0:47]));
ice1f_array_LT_top I_lt_col_t09 ( .glb_netwk_to(net1310[0:7]),
     .glb_netwk_bo(net1424[0:7]), .vdd_cntl(vdd_cntl_r[127:0]),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .top_op_08({slf_op_23_17[3], slf_op_23_17[2], slf_op_23_17[1],
     slf_op_23_17[0], slf_op_23_17[3], slf_op_23_17[2],
     slf_op_23_17[1], slf_op_23_17[0]}), .tnl_op_08({slf_op_22_17[3],
     slf_op_22_17[2], slf_op_22_17[1], slf_op_22_17[0],
     slf_op_22_17[3], slf_op_22_17[2], slf_op_22_17[1],
     slf_op_22_17[0]}), .tnr_op_08({slf_op_12_17[3], slf_op_12_17[2],
     slf_op_12_17[1], slf_op_12_17[0], slf_op_12_17[3],
     slf_op_12_17[2], slf_op_12_17[1], slf_op_12_17[0]}),
     .sp12_v_t_08(net1318[0:23]), .sp4_v_t_08(net1319[0:47]),
     .wl(wl_r[127:0]), .rgt_op_03(net1321[0:7]),
     .slf_op_02(net951[0:7]), .rgt_op_02(net1323[0:7]),
     .rgt_op_01(slf_op_10_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net1145[0:7]), .lft_op_03(net1135[0:7]),
     .lft_op_02(net1137[0:7]), .lft_op_01(slf_op_08_09[7:0]),
     .rgt_op_04(net1331[0:7]), .carry_in(carry_in_09_09),
     .bnl_op_01(bnl_op_09_09[7:0]), .slf_op_04(net959[0:7]),
     .slf_op_03(net949[0:7]), .slf_op_01(slf_op_09_09[7:0]),
     .sp4_h_l_04(net978[0:47]), .carry_out(net1434),
     .sp12_v_b__01(sp12_v_b_09_09[23:0]), .sp12_h_r_04(net1340[0:23]),
     .sp12_h_r_03(net1341[0:23]), .sp12_h_r_02(net1342[0:23]),
     .sp12_h_r_01(net1343[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_09_09[47:0]), .sp4_r_v_b_04(net1346[0:47]),
     .sp4_r_v_b_03(net1347[0:47]), .sp4_r_v_b_02(net1348[0:47]),
     .sp4_r_v_b_01(sp4_v_b_10_09[47:0]), .sp4_h_r_04(net1350[0:47]),
     .sp4_h_r_03(net1351[0:47]), .sp4_h_r_02(net1352[0:47]),
     .sp4_h_r_01(net1353[0:47]), .sp4_h_l_03(net979[0:47]),
     .sp4_h_l_02(net980[0:47]), .sp4_h_l_01(net981[0:47]),
     .bl(bl[161:108]), .bot_op_01(bot_op_09_09[7:0]),
     .sp12_h_l_01(net971[0:23]), .sp12_h_l_02(net970[0:23]),
     .sp12_h_l_03(net969[0:23]), .sp12_h_l_04(net968[0:23]),
     .sp4_v_b_04(net974[0:47]), .sp4_v_b_03(net975[0:47]),
     .sp4_v_b_02(net976[0:47]), .bnr_op_01(bnr_op_09_09[7:0]),
     .sp4_h_l_05(net1002[0:47]), .sp4_h_l_06(net1001[0:47]),
     .sp4_h_l_07(net1000[0:47]), .sp4_h_l_08(net999[0:47]),
     .sp4_h_r_08(net1371[0:47]), .sp4_h_r_07(net1372[0:47]),
     .sp4_h_r_06(net1373[0:47]), .sp4_h_r_05(net1374[0:47]),
     .slf_op_05(net1010[0:7]), .slf_op_06(net1009[0:7]),
     .slf_op_07(net1008[0:7]), .slf_op_08(net1438[0:7]),
     .rgt_op_08(net1441[0:7]), .rgt_op_07(net1380[0:7]),
     .rgt_op_06(net1381[0:7]), .rgt_op_05(net1382[0:7]),
     .lft_op_08(net1430[0:7]), .lft_op_07(net1194[0:7]),
     .lft_op_06(net1195[0:7]), .lft_op_05(net1196[0:7]),
     .sp12_h_l_08(net1021[0:23]), .sp12_h_l_07(net1020[0:23]),
     .sp12_h_l_06(net1019[0:23]), .sp12_h_r_05(net1390[0:23]),
     .sp12_h_r_06(net1391[0:23]), .sp12_h_r_07(net1392[0:23]),
     .sp12_h_r_08(net1393[0:23]), .sp12_h_l_05(net1018[0:23]),
     .sp4_r_v_b_05(net1395[0:47]), .sp4_r_v_b_06(net1396[0:47]),
     .sp4_r_v_b_07(net1397[0:47]), .sp4_r_v_b_08(net1398[0:47]),
     .sp4_v_b_08(net1026[0:47]), .sp4_v_b_07(net1025[0:47]),
     .sp4_v_b_06(net1024[0:47]), .sp4_v_b_05(net1023[0:47]));
fabric_outbuf12p I_fbuf_f1310 ( .fabric_out(net_fabric_out_13_10),
     .cout(fabric_out_13_10));
fabric_outbuf12p I_fbuf_f0817 ( .fabric_out(net_fabric_out_08_17),
     .cout(fabric_out_08_17));
fabric_outbuf12p I_fbuf_p0717a ( .fabric_out(padinlat_t_r[0]),
     .cout(padin_07_17a));
fabric_outbuf12p I_fbuf_f0717 ( .fabric_out(net_fabric_out_07_17),
     .cout(fabric_out_07_17));
fabric_outbuf12p I_fbuf_p1309a ( .fabric_out(padinlat_r[0]),
     .cout(padin_13_09a));
fabric_outbuf12p I_fbuf_f1309 ( .fabric_out(net_fabric_out_13_09),
     .cout(fabric_out_13_09));
clk_quad_buf12px8 I_clk_quad_buf12px8_tr ( .clko(clk_tree_drv[7:0]),
     .clki(glb_in[7:0]));

endmodule
// Library - leafcell, Cell - ice1f_array_LFT_IO_top12io, View -
//schematic
// LAST TIME SAVED: Jul 17 09:08:37 2009
// NETLIST TIME: Aug 24 09:59:02 2009
`timescale 1ns / 1ns 

module ice1f_array_LFT_IO_top12io ( cf_l, fabric_out_09, fabric_out_10,
     fabric_out_11, fabric_out_12, fabric_out_13, fabric_out_14,
     fabric_out_15, fabric_out_16, padeb, pado, sdo, slf_op_00_09,
     slf_op_00_10, slf_op_00_11, slf_op_00_12, slf_op_00_13,
     slf_op_00_14, slf_op_00_15, slf_op_00_16, spi_ss_in_b,
     SP4_h_l_00_09, SP4_h_l_00_10, SP4_h_l_00_11, SP4_h_l_00_12,
     SP4_h_l_00_13, SP4_h_l_00_14, SP4_h_l_00_15, SP4_h_l_00_16,
     SP12_h_l_00_09, SP12_h_l_00_10, SP12_h_l_00_11, SP12_h_l_00_12,
     SP12_h_l_00_13, SP12_h_l_00_14, SP12_h_l_00_15, SP12_h_l_00_16,
     bl, pgate, reset_b, sp4_v_b_00_16, sp4_v_t_00_09, vdd_cntl, wl,
     bnl_op_00_09, bs_en, cdone_in, ceb, glb_netwk_col, hiz_b, hold,
     mode, padin, prog, r, rgt_op_00_09, rgt_op_00_10, rgt_op_00_11,
     rgt_op_00_12, rgt_op_00_13, rgt_op_00_14, rgt_op_00_15,
     rgt_op_00_16, sdi, shift, spioeb, spiout, tclk, tnr_op_00_09,
     update );
output  fabric_out_09, fabric_out_10, fabric_out_11, fabric_out_12,
     fabric_out_13, fabric_out_14, fabric_out_15, fabric_out_16, sdo;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_00_11;
output [3:0]  slf_op_00_13;
output [3:0]  slf_op_00_10;
output [3:0]  slf_op_00_15;
output [3:0]  slf_op_00_16;
output [3:0]  slf_op_00_09;
output [3:0]  slf_op_00_12;
output [3:0]  slf_op_00_14;
output [11:0]  pado;
output [11:0]  padeb;
output [191:0]  cf_l;
output [15:0]  spi_ss_in_b;

inout [23:0]  SP12_h_l_00_10;
inout [47:0]  SP4_h_l_00_16;
inout [47:0]  SP4_h_l_00_14;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_00_12;
inout [23:0]  SP12_h_l_00_09;
inout [15:0]  sp4_v_b_00_16;
inout [23:0]  SP12_h_l_00_14;
inout [23:0]  SP12_h_l_00_11;
inout [23:0]  SP12_h_l_00_13;
inout [47:0]  SP4_h_l_00_15;
inout [15:0]  sp4_v_t_00_09;
inout [23:0]  SP12_h_l_00_15;
inout [47:0]  SP4_h_l_00_10;
inout [23:0]  SP12_h_l_00_16;
inout [47:0]  SP4_h_l_00_11;
inout [47:0]  SP4_h_l_00_13;
inout [127:0]  vdd_cntl;
inout [127:0]  reset_b;
inout [47:0]  SP4_h_l_00_09;
inout [23:0]  SP12_h_l_00_12;
inout [127:0]  pgate;
inout [127:0]  wl;

input [7:0]  rgt_op_00_14;
input [7:0]  rgt_op_00_11;
input [7:0]  rgt_op_00_13;
input [7:0]  rgt_op_00_12;
input [7:0]  rgt_op_00_09;
input [7:0]  bnl_op_00_09;
input [7:0]  rgt_op_00_15;
input [7:0]  glb_netwk_col;
input [16:9]  cdone_in;
input [7:0]  rgt_op_00_16;
input [11:0]  padin;
input [7:0]  tnr_op_00_09;
input [15:0]  spiout;
input [15:0]  spioeb;
input [7:0]  rgt_op_00_10;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net348;

wire  [0:15]  net385;

wire  [1:0]  noconn0015;

wire  [7:0]  colbuf_cntl_b;

wire  [0:7]  net621;

wire  [0:15]  net529;

wire  [0:7]  net622;

wire  [0:7]  net628;

wire  [7:0]  glb_netwk_t;

wire  [0:15]  net601;

wire  [0:15]  net421;

wire  [0:1]  net384;

wire  [0:15]  net493;

wire  [0:7]  net512;

wire  [7:0]  colbuf_cntl_t;

wire  [0:15]  net457;

wire  [0:7]  net638;

wire  [0:1]  net347;

wire  [7:0]  glb_netwk_b;

wire  [0:15]  net565;

wire  [0:7]  net629;



clk_colbuf1kx8 I_clk_colbuf1kx8_t ( .colbuf_cntl(colbuf_cntl_t[7:0]),
     .col_clk(glb_netwk_t[7:0]), .clk_in(glb_netwk_col[7:0]));
clk_colbuf1kx8 I_clk_colbuf1kx8_b ( .colbuf_cntl(colbuf_cntl_b[7:0]),
     .col_clk(glb_netwk_b[7:0]), .clk_in(glb_netwk_col[7:0]));
io_col4_LFT_rev I_io_00_16 ( .cbit_colcntl(net621[0:7]), .ceb(ceb),
     .sdo(net371), .sdi(sdi), .spiout(spiout[15:14]),
     .cdone_in(cdone_in[16]), .spioeb(spioeb[15:14]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(net347[0:1]), .pado(net347[0:1]),
     .padeb(net348[0:1]), .sp4_v_t(sp4_v_t_00_09[15:0]),
     .sp4_h_l(SP4_h_l_00_16[47:0]), .sp12_h_l(SP12_h_l_00_16[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[15:14]),
     .tnl_op(tnr_op_00_09[7:0]), .lft_op(rgt_op_00_16[7:0]),
     .bnl_op(rgt_op_00_15[7:0]), .pgate(pgate[127:112]),
     .reset(reset_b[127:112]), .sp4_v_b(net385[0:15]),
     .wl(wl[127:112]), .cf(cf_l[191:168]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[127:112]), .slf_op(slf_op_00_16[3:0]),
     .glb_netwk(glb_netwk_t[7:0]), .hold(hold),
     .fabric_out(fabric_out_16));
io_col4_LFT_rev I_io_00_15 ( .cbit_colcntl(net622[0:7]), .ceb(ceb),
     .sdo(net443), .sdi(net371), .spiout(spiout[13:12]),
     .cdone_in(cdone_in[15]), .spioeb(spioeb[13:12]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(noconn0015[1:0]), .pado(noconn0015[1:0]),
     .padeb(net384[0:1]), .sp4_v_t(net385[0:15]),
     .sp4_h_l(SP4_h_l_00_15[47:0]), .sp12_h_l(SP12_h_l_00_15[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[13:12]),
     .tnl_op(rgt_op_00_16[7:0]), .lft_op(rgt_op_00_15[7:0]),
     .bnl_op(rgt_op_00_14[7:0]), .pgate(pgate[111:96]),
     .reset(reset_b[111:96]), .sp4_v_b(net457[0:15]), .wl(wl[111:96]),
     .cf(cf_l[167:144]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_00_15[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_15));
io_col4_LFT_rev I_io_00_13 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net587), .sdi(net407), .spiout(spiout[9:8]),
     .cdone_in(cdone_in[13]), .spioeb(spioeb[9:8]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[9:8]), .pado(pado[9:8]),
     .padeb(padeb[9:8]), .sp4_v_t(net421[0:15]),
     .sp4_h_l(SP4_h_l_00_13[47:0]), .sp12_h_l(SP12_h_l_00_13[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[9:8]),
     .tnl_op(rgt_op_00_14[7:0]), .lft_op(rgt_op_00_13[7:0]),
     .bnl_op(rgt_op_00_12[7:0]), .pgate(pgate[79:64]),
     .reset(reset_b[79:64]), .sp4_v_b(net601[0:15]), .wl(wl[79:64]),
     .cf(cf_l[119:96]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_00_13[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_13));
io_col4_LFT_rev I_io_00_14 ( .cbit_colcntl(net638[0:7]), .ceb(ceb),
     .sdo(net407), .sdi(net443), .spiout(spiout[11:10]),
     .cdone_in(cdone_in[14]), .spioeb(spioeb[11:10]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[11:10]), .pado(pado[11:10]),
     .padeb(padeb[11:10]), .sp4_v_t(net457[0:15]),
     .sp4_h_l(SP4_h_l_00_14[47:0]), .sp12_h_l(SP12_h_l_00_14[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[11:10]),
     .tnl_op(rgt_op_00_15[7:0]), .lft_op(rgt_op_00_14[7:0]),
     .bnl_op(rgt_op_00_13[7:0]), .pgate(pgate[95:80]),
     .reset(reset_b[95:80]), .sp4_v_b(net421[0:15]), .wl(wl[95:80]),
     .cf(cf_l[143:120]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_00_14[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_14));
io_col4_LFT_rev I_io_00_10 ( .cbit_colcntl(net628[0:7]), .ceb(ceb),
     .sdo(net515), .sdi(net479), .spiout(spiout[3:2]),
     .cdone_in(cdone_in[10]), .spioeb(spioeb[3:2]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[3:2]), .pado(pado[3:2]),
     .padeb(padeb[3:2]), .sp4_v_t(net493[0:15]),
     .sp4_h_l(SP4_h_l_00_10[47:0]), .sp12_h_l(SP12_h_l_00_10[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[3:2]),
     .tnl_op(rgt_op_00_11[7:0]), .lft_op(rgt_op_00_10[7:0]),
     .bnl_op(rgt_op_00_09[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b(net529[0:15]), .wl(wl[31:16]),
     .cf(cf_l[47:24]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_00_10[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_10));
io_col4_LFT_rev I_io_00_09 ( .cbit_colcntl(net512[0:7]), .ceb(ceb),
     .sdo(sdo), .sdi(net515), .spiout(spiout[1:0]),
     .cdone_in(cdone_in[9]), .spioeb(spioeb[1:0]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .sp4_v_t(net529[0:15]),
     .sp4_h_l(SP4_h_l_00_09[47:0]), .sp12_h_l(SP12_h_l_00_09[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[1:0]),
     .tnl_op(rgt_op_00_10[7:0]), .lft_op(rgt_op_00_09[7:0]),
     .bnl_op(bnl_op_00_09[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(sp4_v_b_00_16[15:0]),
     .wl(wl[15:0]), .cf(cf_l[23:0]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_00_09[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold),
     .fabric_out(fabric_out_09));
io_col4_LFT_rev I_io_00_11 ( .cbit_colcntl(net629[0:7]), .ceb(ceb),
     .sdo(net479), .sdi(net551), .spiout(spiout[5:4]),
     .cdone_in(cdone_in[11]), .spioeb(spioeb[5:4]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[5:4]), .pado(pado[5:4]),
     .padeb(padeb[5:4]), .sp4_v_t(net565[0:15]),
     .sp4_h_l(SP4_h_l_00_11[47:0]), .sp12_h_l(SP12_h_l_00_11[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[5:4]),
     .tnl_op(rgt_op_00_12[7:0]), .lft_op(rgt_op_00_11[7:0]),
     .bnl_op(rgt_op_00_10[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b(net493[0:15]), .wl(wl[47:32]),
     .cf(cf_l[71:48]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_00_11[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_11));
io_col4_LFT_rev I_io_00_12 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net551), .sdi(net587), .spiout(spiout[7:6]),
     .cdone_in(cdone_in[12]), .spioeb(spioeb[7:6]), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk),
     .update(update), .padin(padin[7:6]), .pado(pado[7:6]),
     .padeb(padeb[7:6]), .sp4_v_t(net601[0:15]),
     .sp4_h_l(SP4_h_l_00_12[47:0]), .sp12_h_l(SP12_h_l_00_12[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[7:6]),
     .tnl_op(rgt_op_00_13[7:0]), .lft_op(rgt_op_00_12[7:0]),
     .bnl_op(rgt_op_00_11[7:0]), .pgate(pgate[63:48]),
     .reset(reset_b[63:48]), .sp4_v_b(net565[0:15]), .wl(wl[63:48]),
     .cf(cf_l[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_00_12[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_12));

endmodule
// Library - leafcell, Cell - ice1f_array_TOP_IO_lft, View - schematic
// LAST TIME SAVED: Jun 30 15:10:18 2009
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module ice1f_array_TOP_IO_lft ( bs_en_o, ceb_o, cf_top_l,
     fabric_out_06_17, hiz_b_o, mode_o, padeb_t_l, pado_t_l, r_o, sdo,
     shift_o, slf_op_01_17, slf_op_02_17, slf_op_03_17, slf_op_04_17,
     slf_op_05_17, slf_op_06_17, tclk_o, update_o, bl_01, bl_02, bl_03,
     bl_04, bl_05, bl_06, sp4_h_l_01_17, sp4_h_r_06_17, sp4_v_b_01_17,
     sp4_v_b_02_17, sp4_v_b_03_17, sp4_v_b_04_17, sp4_v_b_05_17,
     sp4_v_b_06_17, sp12_v_b_01_17, sp12_v_b_02_17, sp12_v_b_03_17,
     sp12_v_b_04_17, sp12_v_b_05_17, sp12_v_b_06_17, bnl_op_01_17,
     bnr_op_06_17, bs_en_i, ceb_i, end_of_startup_top_l, glb_net_01,
     glb_net_02, glb_net_03, glb_net_04, glb_net_05, glb_net_06,
     hiz_b_i, hold_t_l, lft_op_01_17, lft_op_02_17, lft_op_03_17,
     lft_op_04_17, lft_op_05_17, lft_op_06_17, mode_i, padin_t_l,
     pgate_l, prog, r_i, reset_l, sdi, shift_i, tclk_i, tiegnd, tievdd,
     update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_06_17, hiz_b_o, mode_o, r_o, sdo,
     shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, tiegnd, tievdd, update_i;

output [3:0]  slf_op_06_17;
output [3:0]  slf_op_04_17;
output [3:0]  slf_op_05_17;
output [3:0]  slf_op_01_17;
output [11:0]  padeb_t_l;
output [3:0]  slf_op_03_17;
output [3:0]  slf_op_02_17;
output [143:0]  cf_top_l;
output [11:0]  pado_t_l;

inout [47:0]  sp4_v_b_02_17;
inout [47:0]  sp4_v_b_04_17;
inout [23:0]  sp12_v_b_01_17;
inout [47:0]  sp4_v_b_05_17;
inout [23:0]  sp12_v_b_05_17;
inout [47:0]  sp4_v_b_01_17;
inout [15:0]  sp4_h_l_01_17;
inout [23:0]  sp12_v_b_04_17;
inout [23:0]  sp12_v_b_03_17;
inout [47:0]  sp4_v_b_06_17;
inout [53:0]  bl_04;
inout [23:0]  sp12_v_b_06_17;
inout [53:0]  bl_01;
inout [53:0]  bl_05;
inout [15:0]  sp4_h_r_06_17;
inout [53:0]  bl_02;
inout [47:0]  sp4_v_b_03_17;
inout [41:0]  bl_03;
inout [23:0]  sp12_v_b_02_17;
inout [53:0]  bl_06;

input [15:0]  vdd_cntl_l;
input [7:0]  lft_op_03_17;
input [15:0]  reset_l;
input [7:0]  bnr_op_06_17;
input [7:0]  glb_net_01;
input [7:0]  glb_net_06;
input [7:0]  glb_net_04;
input [15:0]  wl_l;
input [15:0]  pgate_l;
input [7:0]  bnl_op_01_17;
input [7:0]  lft_op_04_17;
input [7:0]  glb_net_05;
input [7:0]  glb_net_02;
input [7:0]  lft_op_05_17;
input [7:0]  glb_net_03;
input [7:0]  lft_op_06_17;
input [7:0]  lft_op_02_17;
input [7:0]  lft_op_01_17;
input [6:1]  end_of_startup_top_l;
input [11:0]  padin_t_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net533;

wire  [0:15]  net369;

wire  [0:1]  net547;

wire  [0:1]  net373;

wire  [0:1]  net538;

wire  [0:1]  net543;

wire  [0:1]  net544;

wire  [0:15]  net334;

wire  [0:15]  net439;

wire  [0:15]  net474;

wire  [0:15]  net404;



io_col4_TOP_rev I_io_t01 ( .sdo(net303), .sdi(net319), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[1]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_01_17[15:0]), .mode(mode_i),
     .shift(shift_i), .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i),
     .tclk(tclk_i), .update(update_i), .padin(padin_t_l[1:0]),
     .pado(pado_t_l[1:0]), .padeb(padeb_t_l[1:0]),
     .sp4_v_b(net334[0:15]), .sp4_h_l(sp4_v_b_01_17[47:0]),
     .sp12_h_l(sp12_v_b_01_17[23:0]), .prog(prog),
     .spi_ss_in_b(net544[0:1]), .tnl_op(bnl_op_01_17[7:0]),
     .lft_op(lft_op_01_17[7:0]), .bnl_op(lft_op_02_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_01[5],
     bl_01[4], bl_01[37], bl_01[36], bl_01[35], bl_01[34], bl_01[33],
     bl_01[32], bl_01[14], bl_01[20], bl_01[19], bl_01[18], bl_01[17],
     bl_01[16], bl_01[27], bl_01[26], bl_01[25], bl_01[23]}),
     .wl(wl_l[15:0]), .cf(cf_top_l[23:0]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_01_17[3:0]),
     .glb_netwk(glb_net_01[7:0]), .hold(hold_t_l),
     .fabric_out(net534));
io_col4_TOP_rev I_io_t02 ( .sdo(net319), .sdi(net354), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[2]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net334[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_l[3:2]), .pado(pado_t_l[3:2]),
     .padeb(padeb_t_l[3:2]), .sp4_v_b(net369[0:15]),
     .sp4_h_l(sp4_v_b_02_17[47:0]), .sp12_h_l(sp12_v_b_02_17[23:0]),
     .prog(prog), .spi_ss_in_b(net373[0:1]),
     .tnl_op(lft_op_01_17[7:0]), .lft_op(lft_op_02_17[7:0]),
     .bnl_op(lft_op_03_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[47:24]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_17[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_t_l), .fabric_out(net387));
io_col4_TOP_rev I_io_t03 ( .sdo(net354), .sdi(net389), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[3]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net369[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_l[5:4]), .pado(pado_t_l[5:4]),
     .padeb(padeb_t_l[5:4]), .sp4_v_b(net404[0:15]),
     .sp4_h_l(sp4_v_b_03_17[47:0]), .sp12_h_l(sp12_v_b_03_17[23:0]),
     .prog(prog), .spi_ss_in_b(net533[0:1]),
     .tnl_op(lft_op_02_17[7:0]), .lft_op(lft_op_03_17[7:0]),
     .bnl_op(lft_op_04_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[71:48]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_17[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_t_l), .fabric_out(net422));
io_col4_TOP_rev I_io_t05 ( .sdo(net459), .sdi(net424), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[5]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net474[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_l[9:8]), .pado(pado_t_l[9:8]),
     .padeb(padeb_t_l[9:8]), .sp4_v_b(net439[0:15]),
     .sp4_h_l(sp4_v_b_05_17[47:0]), .sp12_h_l(sp12_v_b_05_17[23:0]),
     .prog(prog), .spi_ss_in_b(net538[0:1]),
     .tnl_op(lft_op_04_17[7:0]), .lft_op(lft_op_05_17[7:0]),
     .bnl_op(lft_op_06_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[119:96]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_17[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_t_l), .fabric_out(net539));
io_col4_TOP_rev I_io_t04 ( .sdo(net389), .sdi(net459), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[4]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net404[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_l[7:6]), .pado(pado_t_l[7:6]),
     .padeb(padeb_t_l[7:6]), .sp4_v_b(net474[0:15]),
     .sp4_h_l(sp4_v_b_04_17[47:0]), .sp12_h_l(sp12_v_b_04_17[23:0]),
     .prog(prog), .spi_ss_in_b(net543[0:1]),
     .tnl_op(lft_op_03_17[7:0]), .lft_op(lft_op_04_17[7:0]),
     .bnl_op(lft_op_05_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_04[5], bl_04[4], bl_04[37],
     bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32], bl_04[14],
     bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16], bl_04[27],
     bl_04[26], bl_04[25], bl_04[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[95:72]), .ceb(ceb_i), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_17[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_t_l), .fabric_out(net542));
io_col4_TOP_rev I_io_t06 ( .sdo(net424), .sdi(sdi), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_l[6]), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net439[0:15]), .mode(mode_i), .shift(shift_i),
     .hiz_b(hiz_b_i), .r(r_i), .bs_en(bs_en_i), .tclk(tclk_i),
     .update(update_i), .padin(padin_t_l[11:10]),
     .pado(pado_t_l[11:10]), .padeb(padeb_t_l[11:10]),
     .sp4_v_b(sp4_h_r_06_17[15:0]), .sp4_h_l(sp4_v_b_06_17[47:0]),
     .sp12_h_l(sp12_v_b_06_17[23:0]), .prog(prog),
     .spi_ss_in_b(net547[0:1]), .tnl_op(lft_op_05_17[7:0]),
     .lft_op(lft_op_06_17[7:0]), .bnl_op(bnr_op_06_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_06[5],
     bl_06[4], bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33],
     bl_06[32], bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17],
     bl_06[16], bl_06[27], bl_06[26], bl_06[25], bl_06[23]}),
     .wl(wl_l[15:0]), .cf(cf_top_l[143:120]), .ceb(ceb_i),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_06_17[3:0]),
     .glb_netwk(glb_net_06[7:0]), .hold(hold_t_l),
     .fabric_out(fabric_out_06_17));
scanbuf1f I_scanbuf_tl ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(net303), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(tclk_o), .shift_o(shift_o),
     .sdo(sdo), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));

endmodule
// Library - leafcell, Cell - ice1f_quad_tl, View - schematic
// LAST TIME SAVED: Jul 22 09:24:43 2009
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module ice1f_quad_tl ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, ceb_o, cf_l, cf_t, fabric_out_00_09,
     fabric_out_06_17, hiz_b_o, mode_o, padeb_l_t, padeb_t_l,
     padin_00_09a, padin_06_17b, pado_l_t, pado_t_l, r_o, sdo, shift_o,
     slf_op_00_09, slf_op_01_09, slf_op_02_09, slf_op_03_09,
     slf_op_04_09, slf_op_05_09, slf_op_06_09, slf_op_06_10,
     slf_op_06_11, slf_op_06_12, slf_op_06_13, slf_op_06_14,
     slf_op_06_15, slf_op_06_16, slf_op_06_17, tclk_o, update_o, bl,
     pgate_l, reset_b_l, sp4_h_r_06_09, sp4_h_r_06_10, sp4_h_r_06_11,
     sp4_h_r_06_12, sp4_h_r_06_13, sp4_h_r_06_14, sp4_h_r_06_15,
     sp4_h_r_06_16, sp4_h_r_06_17, sp4_r_v_b_06_09, sp4_r_v_b_06_10,
     sp4_r_v_b_06_11, sp4_r_v_b_06_12, sp4_r_v_b_06_13,
     sp4_r_v_b_06_14, sp4_r_v_b_06_15, sp4_r_v_b_06_16, sp4_v_b_00_09,
     sp4_v_b_01_09, sp4_v_b_02_09, sp4_v_b_03_09, sp4_v_b_04_09,
     sp4_v_b_05_09, sp4_v_b_06_09, sp12_h_r_06_09, sp12_h_r_06_10,
     sp12_h_r_06_11, sp12_h_r_06_12, sp12_h_r_06_13, sp12_h_r_06_14,
     sp12_h_r_06_15, sp12_h_r_06_16, sp12_v_b_01_09, sp12_v_b_02_09,
     sp12_v_b_03_09, sp12_v_b_04_09, sp12_v_b_05_09, sp12_v_b_06_09,
     vdd_cntl_l, wl_l, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_01_09, bnl_op_02_09, bnl_op_03_09,
     bnl_op_04_09, bnl_op_05_09, bnl_op_06_09, bnr_op_00_09,
     bnr_op_01_09, bnr_op_02_09, bnr_op_03_09, bnr_op_04_09,
     bnr_op_05_09, bnr_op_06_09, bot_op_01_09, bot_op_02_09,
     bot_op_03_09, bot_op_04_09, bot_op_05_09, bot_op_06_09, bs_en_i,
     carry_in_01_09, carry_in_02_09, carry_in_04_09, carry_in_05_09,
     carry_in_06_09, ceb_i, end_of_startup_lft_t, end_of_startup_top_l,
     glb_in, hiz_b_i, hold_l_t, hold_t_l, last_rsr, mode_i, padin_l_t,
     padin_t_l, prog, purst, r_i, rgt_op_06_09, rgt_op_06_10,
     rgt_op_06_11, rgt_op_06_12, rgt_op_06_13, rgt_op_06_14,
     rgt_op_06_15, rgt_op_06_16, sdi, shift_i, tclk_i, tiegnd, tievdd,
     tnr_op_06_16, update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bs_en_o, ceb_o,
     fabric_out_00_09, fabric_out_06_17, hiz_b_o, mode_o, padin_00_09a,
     padin_06_17b, r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en_i,
     carry_in_01_09, carry_in_02_09, carry_in_04_09, carry_in_05_09,
     carry_in_06_09, ceb_i, hiz_b_i, hold_l_t, hold_t_l, last_rsr,
     mode_i, prog, purst, r_i, sdi, shift_i, tclk_i, tiegnd, tievdd,
     update_i;

output [7:0]  slf_op_06_11;
output [11:0]  pado_l_t;
output [7:0]  slf_op_06_13;
output [7:0]  slf_op_06_12;
output [7:0]  slf_op_01_09;
output [7:0]  slf_op_02_09;
output [11:0]  padeb_t_l;
output [7:0]  slf_op_06_15;
output [7:0]  bm_sa_o;
output [11:0]  padeb_l_t;
output [7:0]  slf_op_06_10;
output [7:0]  slf_op_05_09;
output [7:0]  slf_op_04_09;
output [143:0]  cf_t;
output [7:0]  slf_op_06_09;
output [191:0]  cf_l;
output [3:0]  slf_op_06_17;
output [11:0]  pado_t_l;
output [3:0]  slf_op_00_09;
output [7:0]  slf_op_06_16;
output [7:0]  slf_op_03_09;
output [7:0]  slf_op_06_14;

inout [23:0]  sp12_h_r_06_14;
inout [47:0]  sp4_h_r_06_14;
inout [47:0]  sp4_h_r_06_15;
inout [23:0]  sp12_h_r_06_12;
inout [47:0]  sp4_r_v_b_06_09;
inout [47:0]  sp4_r_v_b_06_11;
inout [47:0]  sp4_h_r_06_16;
inout [23:0]  sp12_h_r_06_11;
inout [23:0]  sp12_h_r_06_10;
inout [47:0]  sp4_r_v_b_06_13;
inout [23:0]  sp12_v_b_01_09;
inout [143:0]  reset_b_l;
inout [47:0]  sp4_r_v_b_06_12;
inout [47:0]  sp4_v_b_02_09;
inout [15:0]  sp4_h_r_06_17;
inout [15:0]  sp4_v_b_00_09;
inout [23:0]  sp12_v_b_04_09;
inout [47:0]  sp4_v_b_03_09;
inout [47:0]  sp4_v_b_04_09;
inout [47:0]  sp4_r_v_b_06_14;
inout [23:0]  sp12_h_r_06_15;
inout [47:0]  sp4_h_r_06_12;
inout [47:0]  sp4_v_b_05_09;
inout [23:0]  sp12_v_b_03_09;
inout [47:0]  sp4_h_r_06_11;
inout [143:0]  pgate_l;
inout [47:0]  sp4_r_v_b_06_10;
inout [47:0]  sp4_v_b_01_09;
inout [47:0]  sp4_h_r_06_09;
inout [47:0]  sp4_r_v_b_06_15;
inout [47:0]  sp4_h_r_06_13;
inout [23:0]  sp12_v_b_02_09;
inout [47:0]  sp4_v_b_06_09;
inout [143:0]  vdd_cntl_l;
inout [23:0]  sp12_v_b_05_09;
inout [329:0]  bl;
inout [23:0]  sp12_h_r_06_09;
inout [23:0]  sp12_h_r_06_13;
inout [143:0]  wl_l;
inout [23:0]  sp12_h_r_06_16;
inout [47:0]  sp4_h_r_06_10;
inout [47:0]  sp4_r_v_b_06_16;
inout [23:0]  sp12_v_b_06_09;

input [7:0]  rgt_op_06_09;
input [7:0]  bnl_op_01_09;
input [7:0]  rgt_op_06_15;
input [7:0]  rgt_op_06_13;
input [7:0]  bm_sa_i;
input [7:0]  bot_op_06_09;
input [7:0]  bot_op_03_09;
input [7:0]  bnl_op_03_09;
input [7:0]  bnl_op_04_09;
input [7:0]  bnr_op_01_09;
input [7:0]  bnr_op_03_09;
input [11:0]  padin_l_t;
input [7:0]  bnr_op_06_09;
input [7:0]  bnl_op_05_09;
input [7:0]  rgt_op_06_12;
input [7:0]  bot_op_04_09;
input [7:0]  bnl_op_02_09;
input [7:0]  bot_op_05_09;
input [7:0]  bnr_op_02_09;
input [7:0]  rgt_op_06_10;
input [7:0]  bnr_op_05_09;
input [7:0]  rgt_op_06_16;
input [7:0]  bnl_op_06_09;
input [6:1]  end_of_startup_top_l;
input [7:0]  rgt_op_06_11;
input [16:9]  end_of_startup_lft_t;
input [7:0]  bnr_op_00_09;
input [11:0]  padin_t_l;
input [7:0]  rgt_op_06_14;
input [7:0]  glb_in;
input [7:0]  bnr_op_04_09;
input [7:0]  bot_op_01_09;
input [7:0]  bot_op_02_09;
input [3:0]  tnr_op_06_16;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:47]  net1441;

wire  [0:47]  net692;

wire  [0:47]  net1152;

wire  [0:47]  net1362;

wire  [0:7]  net999;

wire  [0:23]  net685;

wire  [0:23]  net1287;

wire  [0:47]  net966;

wire  [0:47]  net879;

wire  [0:47]  net1177;

wire  [0:47]  net1337;

wire  [0:7]  net895;

wire  [0:23]  net1029;

wire  [0:47]  net880;

wire  [0:47]  net1295;

wire  [0:47]  net1292;

wire  [0:47]  net1200;

wire  [0:23]  net1009;

wire  [0:23]  net1383;

wire  [0:47]  net860;

wire  [0:47]  net819;

wire  [0:7]  net1408;

wire  [0:7]  net1445;

wire  [0:47]  net1386;

wire  [0:47]  net1216;

wire  [0:7]  net1300;

wire  [0:23]  net1144;

wire  [0:7]  net823;

wire  [0:7]  net1207;

wire  [0:23]  net1444;

wire  [0:47]  net937;

wire  [0:47]  net1243;

wire  [0:47]  net1435;

wire  [0:7]  net1427;

wire  [3:0]  slf_op_00_16;

wire  [0:47]  net1175;

wire  [0:23]  net1382;

wire  [0:7]  net1410;

wire  [0:7]  net941;

wire  [0:47]  net684;

wire  [0:23]  net1424;

wire  [0:23]  net681;

wire  [0:47]  net989;

wire  [0:23]  net1197;

wire  [0:47]  net1309;

wire  [0:47]  net1016;

wire  [0:23]  net1146;

wire  [0:23]  net959;

wire  [0:47]  net1361;

wire  [0:47]  net919;

wire  [0:47]  net1015;

wire  [0:7]  net1184;

wire  [0:47]  net909;

wire  [0:23]  net960;

wire  [0:7]  net1426;

wire  [0:47]  net1419;

wire  [0:7]  net679;

wire  [0:47]  net1413;

wire  [3:0]  slf_op_04_17;

wire  [0:47]  net664;

wire  [0:47]  net1363;

wire  [0:47]  net1341;

wire  [0:47]  net668;

wire  [0:23]  net1196;

wire  [0:23]  net844;

wire  [0:23]  net821;

wire  [0:47]  net1014;

wire  [0:47]  net1293;

wire  [0:23]  net1289;

wire  [0:23]  net885;

wire  [0:7]  net906;

wire  [0:23]  net1290;

wire  [0:23]  net1380;

wire  [0:47]  net1201;

wire  [0:23]  net843;

wire  [0:47]  net964;

wire  [0:47]  net1270;

wire  [0:47]  net911;

wire  [0:47]  net917;

wire  [0:7]  net1278;

wire  [0:47]  net1388;

wire  [0:23]  net1239;

wire  [0:23]  net1147;

wire  [0:23]  net883;

wire  [0:47]  net1460;

wire  [0:23]  net842;

wire  [0:47]  net1249;

wire  [0:23]  net1332;

wire  [0:7]  net1218;

wire  [0:7]  net1405;

wire  [0:7]  net928;

wire  [0:47]  net1030;

wire  [0:47]  net1475;

wire  [11:11]  padinlat_t_l;

wire  [0:15]  net653;

wire  [0:7]  net900;

wire  [0:47]  net912;

wire  [0:47]  net680;

wire  [0:23]  net1011;

wire  [3:0]  slf_op_00_12;

wire  [0:23]  net669;

wire  [0:47]  net1199;

wire  [0:7]  net998;

wire  [0:47]  net992;

wire  [0:23]  net847;

wire  [0:47]  net1343;

wire  [0:47]  net676;

wire  [0:7]  net897;

wire  [0:7]  net939;

wire  [0:47]  net1340;

wire  [0:23]  net1194;

wire  [0:23]  net1288;

wire  [3:0]  slf_op_00_13;

wire  [0:47]  net1150;

wire  [0:47]  net1176;

wire  [0:47]  net969;

wire  [0:7]  net1127;

wire  [0:23]  net1122;

wire  [0:7]  net898;

wire  [0:47]  net1294;

wire  [0:7]  net1186;

wire  [0:7]  net1021;

wire  [0:7]  net949;

wire  [0:7]  net1114;

wire  [3:0]  slf_op_00_11;

wire  [0:47]  net1157;

wire  [0:23]  net665;

wire  [0:23]  net1330;

wire  [0:23]  net1195;

wire  [0:7]  net1125;

wire  [0:47]  net1385;

wire  [0:7]  net1022;

wire  [0:23]  net840;

wire  [0:23]  net673;

wire  [3:0]  slf_op_05_17;

wire  [0:7]  net675;

wire  [0:7]  net683;

wire  [0:23]  net1381;

wire  [0:47]  net858;

wire  [0:47]  net1268;

wire  [0:7]  net1406;

wire  [0:47]  net910;

wire  [0:47]  net965;

wire  [0:47]  net971;

wire  [3:0]  slf_op_00_15;

wire  [0:23]  net887;

wire  [0:47]  net1412;

wire  [0:7]  net695;

wire  [0:47]  net1271;

wire  [0:23]  net1238;

wire  [0:23]  net1333;

wire  [0:47]  net1156;

wire  [0:47]  net856;

wire  [0:47]  net1248;

wire  [0:23]  net936;

wire  [3:0]  slf_op_01_17;

wire  [0:7]  net1220;

wire  [0:47]  net1336;

wire  [0:23]  net1008;

wire  [0:47]  net1387;

wire  [0:47]  net878;

wire  [0:7]  net1135;

wire  [0:47]  net968;

wire  [0:7]  net1185;

wire  [0:47]  net672;

wire  [0:7]  net894;

wire  [0:47]  net1244;

wire  [3:0]  slf_op_02_17;

wire  [0:23]  net1215;

wire  [0:47]  net1155;

wire  [0:23]  net1240;

wire  [0:47]  net1250;

wire  [0:7]  net907;

wire  [0:47]  net881;

wire  [0:47]  net863;

wire  [0:7]  net691;

wire  [0:7]  net671;

wire  [3:0]  slf_op_03_17;

wire  [0:47]  net1154;

wire  [0:47]  net1269;

wire  [0:23]  net1331;

wire  [0:47]  net970;

wire  [0:23]  net958;

wire  [0:47]  net861;

wire  [0:47]  net1013;

wire  [0:23]  net1237;

wire  [0:47]  net1342;

wire  [0:15]  net1455;

wire  [0:7]  net687;

wire  [3:0]  slf_op_00_14;

wire  [0:7]  net1228;

wire  [0:47]  net1202;

wire  [0:47]  net1247;

wire  [0:47]  net1245;

wire  [0:23]  net1308;

wire  [3:0]  slf_op_00_10;

wire  [0:47]  net1338;

wire  [0:47]  net1364;

wire  [0:23]  net961;

wire  [0:47]  net1178;

wire  [0:47]  net990;

wire  [0:7]  net1414;

wire  [0:47]  net1123;

wire  [0:47]  net991;

wire  [0:23]  net677;

wire  [0:23]  net1010;

wire  [0:0]  padinlat_l_t;

wire  [0:7]  net1000;

wire  [0:7]  net1279;

wire  [0:47]  net688;

wire  [7:0]  clk_tree_drv;

wire  [0:7]  net1277;

wire  [0:47]  net1151;

wire  [0:23]  net1145;



ice1f_array_LFT_IO_top12io I_preio_lft_t00 ( .padin(padin_l_t[11:0]),
     .pado(pado_l_t[11:0]), .padeb(padeb_l_t[11:0]),
     .cdone_in(end_of_startup_lft_t[16:9]),
     .tnr_op_00_09({slf_op_01_17[3], slf_op_01_17[2], slf_op_01_17[1],
     slf_op_01_17[0], slf_op_01_17[3], slf_op_01_17[2],
     slf_op_01_17[1], slf_op_01_17[0]}), .sp4_v_t_00_09(net653[0:15]),
     .sp4_v_b_00_16(sp4_v_b_00_09[15:0]), .cf_l(cf_l[191:0]),
     .spi_ss_in_b(net1455[0:15]), .spiout({tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, last_rsr}), .spioeb({tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tiegnd}),
     .wl(wl_l[127:0]), .vdd_cntl(vdd_cntl_l[127:0]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .bnl_op_00_09(bnr_op_00_09[7:0]), .SP4_h_l_00_09(net664[0:47]),
     .SP12_h_l_00_09(net665[0:23]), .slf_op_00_09(slf_op_00_09[3:0]),
     .rgt_op_00_09(slf_op_01_09[7:0]), .SP4_h_l_00_10(net668[0:47]),
     .SP12_h_l_00_10(net669[0:23]), .slf_op_00_10(slf_op_00_10[3:0]),
     .rgt_op_00_10(net671[0:7]), .SP4_h_l_00_11(net672[0:47]),
     .SP12_h_l_00_11(net673[0:23]), .slf_op_00_11(slf_op_00_11[3:0]),
     .rgt_op_00_11(net675[0:7]), .SP4_h_l_00_12(net676[0:47]),
     .SP12_h_l_00_12(net677[0:23]), .slf_op_00_12(slf_op_00_12[3:0]),
     .rgt_op_00_12(net679[0:7]), .SP4_h_l_00_13(net680[0:47]),
     .SP12_h_l_00_13(net681[0:23]), .slf_op_00_13(slf_op_00_13[3:0]),
     .rgt_op_00_13(net683[0:7]), .SP4_h_l_00_14(net684[0:47]),
     .SP12_h_l_00_14(net685[0:23]), .slf_op_00_14(slf_op_00_14[3:0]),
     .rgt_op_00_14(net687[0:7]), .SP4_h_l_00_15(net688[0:47]),
     .SP12_h_l_00_15(net1444[0:23]), .slf_op_00_15(slf_op_00_15[3:0]),
     .rgt_op_00_15(net691[0:7]), .SP4_h_l_00_16(net692[0:47]),
     .SP12_h_l_00_16(net1424[0:23]), .slf_op_00_16(slf_op_00_16[3:0]),
     .rgt_op_00_16(net695[0:7]), .fabric_out_09(net_fabric_out_00_09),
     .fabric_out_10(net1411), .fabric_out_11(net1447),
     .fabric_out_12(net1442), .fabric_out_13(net1431),
     .fabric_out_14(net1422), .fabric_out_15(net702),
     .fabric_out_16(net703), .shift(shift_tl), .bs_en(bs_en_tl),
     .mode(mode_tl), .sdi(sdio_tl), .hiz_b(hiz_b_tl), .prog(prog),
     .hold(hold_l_t), .update(update_tl),
     .glb_netwk_col(clk_tree_drv[7:0]), .r(r_tl), .sdo(net731),
     .bl({bl[0], bl[1], bl[2], bl[3], bl[4], bl[5], bl[6], bl[7],
     bl[8], bl[9], bl[10], bl[11], bl[12], bl[13], bl[14], bl[15],
     bl[16], bl[17]}), .tclk(tclk_tl), .ceb(ceb_tl));
pinlatbuf12p I_pinlatbuf12p ( .pad_in(padin_t_l[11]),
     .icegate(hold_t_l), .cbit(cf_t[135]), .cout(padinlat_t_l[11]),
     .prog(prog));
pinlatbuf12p I_pinlatbuf12p_l ( .pad_in(padin_l_t[0]),
     .icegate(hold_l_t), .cbit(cf_l[15]), .cout(padinlat_l_t[0]),
     .prog(prog));
scanbuf1f I_scanbuf_ml ( .update_i(update_tl), .tclk_i(tclk_tl),
     .shift_i(shift_tl), .sdi(net731), .r_i(r_tl), .mode_i(mode_tl),
     .hiz_b_i(hiz_b_tl), .ceb_i(ceb_tl), .bs_en_i(bs_en_tl),
     .update_o(update_o), .tclk_o(tclk_o), .shift_o(shift_o),
     .sdo(sdo), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
ice1f_array_TOP_IO_lft I_preio_top_l ( .padin_t_l(padin_t_l[11:0]),
     .padeb_t_l(padeb_t_l[11:0]), .pado_t_l(pado_t_l[11:0]),
     .bnr_op_06_17(rgt_op_06_16[7:0]), .cf_top_l(cf_t[143:0]),
     .sp4_h_r_06_17(sp4_h_r_06_17[15:0]), .bl_03(bl[167:126]),
     .sp4_h_l_01_17(net653[0:15]), .bnl_op_01_17({slf_op_00_16[3],
     slf_op_00_16[2], slf_op_00_16[1], slf_op_00_16[0],
     slf_op_00_16[3], slf_op_00_16[2], slf_op_00_16[1],
     slf_op_00_16[0]}), .sp4_v_b_01_17(net1216[0:47]),
     .slf_op_01_17(slf_op_01_17[3:0]), .lft_op_01_17(net695[0:7]),
     .sp12_v_b_01_17(net1215[0:23]), .sp4_v_b_02_17(net937[0:47]),
     .slf_op_02_17(slf_op_02_17[3:0]), .lft_op_02_17(net1427[0:7]),
     .sp12_v_b_02_17(net936[0:23]), .sp4_v_b_03_17(net819[0:47]),
     .slf_op_03_17(slf_op_03_17[3:0]), .lft_op_03_17(net1426[0:7]),
     .sp12_v_b_03_17(net821[0:23]), .sp4_v_b_04_17(net1123[0:47]),
     .slf_op_04_17(slf_op_04_17[3:0]), .lft_op_04_17(net895[0:7]),
     .sp12_v_b_04_17(net1122[0:23]), .sp4_v_b_05_17(net1309[0:47]),
     .slf_op_05_17(slf_op_05_17[3:0]), .lft_op_05_17(net1445[0:7]),
     .sp12_v_b_05_17(net1308[0:23]), .sp4_v_b_06_17(net1030[0:47]),
     .slf_op_06_17(slf_op_06_17[3:0]),
     .lft_op_06_17(slf_op_06_16[7:0]), .sp12_v_b_06_17(net1029[0:23]),
     .end_of_startup_top_l(end_of_startup_top_l[6:1]),
     .fabric_out_06_17(net_fabric_out_06_17), .wl_l({wl_l[142],
     wl_l[143], wl_l[141], wl_l[140], wl_l[138], wl_l[139], wl_l[137],
     wl_l[136], wl_l[134], wl_l[135], wl_l[133], wl_l[132], wl_l[130],
     wl_l[131], wl_l[129], wl_l[128]}), .vdd_cntl_l({vdd_cntl_l[142],
     vdd_cntl_l[143], vdd_cntl_l[141], vdd_cntl_l[140],
     vdd_cntl_l[138], vdd_cntl_l[139], vdd_cntl_l[137],
     vdd_cntl_l[136], vdd_cntl_l[134], vdd_cntl_l[135],
     vdd_cntl_l[133], vdd_cntl_l[132], vdd_cntl_l[130],
     vdd_cntl_l[131], vdd_cntl_l[129], vdd_cntl_l[128]}),
     .update_i(update_i), .tievdd(tievdd), .tiegnd(tiegnd),
     .tclk_i(tclk_i), .shift_i(shift_i), .sdi(sdi),
     .reset_l({reset_b_l[142], reset_b_l[143], reset_b_l[141],
     reset_b_l[140], reset_b_l[138], reset_b_l[139], reset_b_l[137],
     reset_b_l[136], reset_b_l[134], reset_b_l[135], reset_b_l[133],
     reset_b_l[132], reset_b_l[130], reset_b_l[131], reset_b_l[129],
     reset_b_l[128]}), .r_i(r_i), .prog(prog), .pgate_l({pgate_l[142],
     pgate_l[143], pgate_l[141], pgate_l[140], pgate_l[138],
     pgate_l[139], pgate_l[137], pgate_l[136], pgate_l[134],
     pgate_l[135], pgate_l[133], pgate_l[132], pgate_l[130],
     pgate_l[131], pgate_l[129], pgate_l[128]}), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .bs_en_i(bs_en_i), .update_o(update_tl),
     .tclk_o(tclk_tl), .shift_o(shift_tl), .sdo(sdio_tl), .r_o(r_tl),
     .mode_o(mode_tl), .hiz_b_o(hiz_b_tl), .glb_net_06(net1021[0:7]),
     .glb_net_05(net1300[0:7]), .glb_net_04(net1114[0:7]),
     .glb_net_03(net823[0:7]), .glb_net_02(net928[0:7]),
     .glb_net_01(net1207[0:7]), .bs_en_o(bs_en_tl),
     .bl_06(bl[329:276]), .bl_05(bl[275:222]), .bl_04(bl[221:168]),
     .bl_02(bl[125:72]), .bl_01(bl[71:18]), .ceb_o(ceb_tl),
     .hold_t_l(hold_t_l), .ceb_i(ceb_i));
ice1f_array_BRAM_top I_bram_col_t03 ( .tnl_op_08({slf_op_02_17[3],
     slf_op_02_17[2], slf_op_02_17[1], slf_op_02_17[0],
     slf_op_02_17[3], slf_op_02_17[2], slf_op_02_17[1],
     slf_op_02_17[0]}), .sp4_v_t_08(net819[0:47]),
     .top_op_08({slf_op_03_17[3], slf_op_03_17[2], slf_op_03_17[1],
     slf_op_03_17[0], slf_op_03_17[3], slf_op_03_17[2],
     slf_op_03_17[1], slf_op_03_17[0]}), .sp12_v_t_08(net821[0:23]),
     .tnr_op_08({slf_op_04_17[3], slf_op_04_17[2], slf_op_04_17[1],
     slf_op_04_17[0], slf_op_04_17[3], slf_op_04_17[2],
     slf_op_04_17[1], slf_op_04_17[0]}), .glb_netwk_top(net823[0:7]),
     .pgate(pgate_l[127:0]), .vdd_cntl(vdd_cntl_l[127:0]),
     .reset_b(reset_b_l[127:0]), .wl(wl_l[127:0]),
     .glb_netwk_bot(net1410[0:7]), .prog(prog),
     .glb_netwk_col(clk_tree_drv[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .sp12_h_l_07(net1010[0:23]), .sp4_v_b_08(net1016[0:47]),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bnr_op_01(bnr_op_03_09[7:0]), .sp12_h_r_06(net840[0:23]),
     .sp12_h_l_06(net1009[0:23]), .sp12_h_r_05(net842[0:23]),
     .sp12_h_r_08(net843[0:23]), .sp12_h_r_03(net844[0:23]),
     .sp12_h_l_08(net1011[0:23]), .sp12_h_l_05(net1008[0:23]),
     .sp12_h_r_07(net847[0:23]), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_sreb_o(bm_sreb_o), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .sp4_r_v_b_01(sp4_v_b_04_09[47:0]),
     .sp4_v_b_02(net966[0:47]), .sp4_r_v_b_02(net856[0:47]),
     .sp4_v_b_03(net965[0:47]), .sp4_r_v_b_03(net858[0:47]),
     .sp4_v_b_04(net964[0:47]), .sp4_r_v_b_04(net860[0:47]),
     .sp4_r_v_b_06(net861[0:47]), .sp4_v_b_06(net1014[0:47]),
     .sp4_r_v_b_05(net863[0:47]), .sp4_v_b_05(net1013[0:47]),
     .lft_op_08(net1427[0:7]), .lft_op_07(net1277[0:7]),
     .lft_op_06(net1278[0:7]), .lft_op_05(net1279[0:7]),
     .sp4_v_b_07(net1015[0:47]), .sp12_h_l_03(net959[0:23]),
     .sp12_h_l_04(net958[0:23]), .sp12_h_l_02(net960[0:23]),
     .sp12_h_l_01(net961[0:23]), .slf_op_07(net998[0:7]),
     .slf_op_08(net1426[0:7]), .sp4_h_l_07(net990[0:47]),
     .sp4_h_l_08(net989[0:47]), .sp4_h_r_07(net878[0:47]),
     .sp4_h_r_08(net879[0:47]), .sp4_r_v_b_07(net880[0:47]),
     .sp4_r_v_b_08(net881[0:47]), .sp4_v_b_01(sp4_v_b_03_09[47:0]),
     .sp12_h_r_01(net883[0:23]), .bm_sdo_i(bm_sdo_i),
     .sp12_h_r_02(net885[0:23]), .bl(bl[167:126]),
     .sp12_h_r_04(net887[0:23]), .sp12_v_b_01(sp12_v_b_03_09[23:0]),
     .bnl_op_01(bnl_op_03_09[7:0]), .lft_op_01(slf_op_02_09[7:0]),
     .lft_op_02(net1220[0:7]), .lft_op_03(net1218[0:7]),
     .lft_op_04(net1228[0:7]), .rgt_op_07(net894[0:7]),
     .rgt_op_08(net895[0:7]), .bot_op_01(bot_op_03_09[7:0]),
     .rgt_op_03(net897[0:7]), .rgt_op_02(net898[0:7]),
     .rgt_op_01(slf_op_04_09[7:0]), .rgt_op_04(net900[0:7]),
     .slf_op_04(net949[0:7]), .slf_op_03(net939[0:7]),
     .slf_op_02(net941[0:7]), .slf_op_01(slf_op_03_09[7:0]),
     .slf_op_06(net999[0:7]), .rgt_op_05(net906[0:7]),
     .rgt_op_06(net907[0:7]), .slf_op_05(net1000[0:7]),
     .sp4_h_r_04(net909[0:47]), .sp4_h_r_03(net910[0:47]),
     .sp4_h_r_02(net911[0:47]), .sp4_h_r_01(net912[0:47]),
     .sp4_h_l_04(net968[0:47]), .sp4_h_l_03(net969[0:47]),
     .sp4_h_l_02(net970[0:47]), .sp4_h_l_01(net971[0:47]),
     .sp4_h_r_06(net917[0:47]), .sp4_h_l_06(net991[0:47]),
     .sp4_h_r_05(net919[0:47]), .sp4_h_l_05(net992[0:47]),
     .bm_sdo_o(bm_sdo_o), .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_sweb_i(bm_sweb_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sweb_o(bm_sweb_o));
ice1f_array_LT_top I_lt_col_t02 ( .glb_netwk_to(net928[0:7]),
     .glb_netwk_bo(net1408[0:7]), .vdd_cntl(vdd_cntl_l[127:0]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .top_op_08({slf_op_02_17[3], slf_op_02_17[2], slf_op_02_17[1],
     slf_op_02_17[0], slf_op_02_17[3], slf_op_02_17[2],
     slf_op_02_17[1], slf_op_02_17[0]}), .tnl_op_08({slf_op_01_17[3],
     slf_op_01_17[2], slf_op_01_17[1], slf_op_01_17[0],
     slf_op_01_17[3], slf_op_01_17[2], slf_op_01_17[1],
     slf_op_01_17[0]}), .tnr_op_08({slf_op_03_17[3], slf_op_03_17[2],
     slf_op_03_17[1], slf_op_03_17[0], slf_op_03_17[3],
     slf_op_03_17[2], slf_op_03_17[1], slf_op_03_17[0]}),
     .sp12_v_t_08(net936[0:23]), .sp4_v_t_08(net937[0:47]),
     .wl(wl_l[127:0]), .rgt_op_03(net939[0:7]),
     .slf_op_02(net1220[0:7]), .rgt_op_02(net941[0:7]),
     .rgt_op_01(slf_op_03_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net679[0:7]), .lft_op_03(net675[0:7]),
     .lft_op_02(net671[0:7]), .lft_op_01(slf_op_01_09[7:0]),
     .rgt_op_04(net949[0:7]), .carry_in(carry_in_02_09),
     .bnl_op_01(bnl_op_02_09[7:0]), .slf_op_04(net1228[0:7]),
     .slf_op_03(net1218[0:7]), .slf_op_01(slf_op_02_09[7:0]),
     .sp4_h_l_04(net1247[0:47]), .carry_out(net956),
     .sp12_v_b__01(sp12_v_b_02_09[23:0]), .sp12_h_r_04(net958[0:23]),
     .sp12_h_r_03(net959[0:23]), .sp12_h_r_02(net960[0:23]),
     .sp12_h_r_01(net961[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_02_09[47:0]), .sp4_r_v_b_04(net964[0:47]),
     .sp4_r_v_b_03(net965[0:47]), .sp4_r_v_b_02(net966[0:47]),
     .sp4_r_v_b_01(sp4_v_b_03_09[47:0]), .sp4_h_r_04(net968[0:47]),
     .sp4_h_r_03(net969[0:47]), .sp4_h_r_02(net970[0:47]),
     .sp4_h_r_01(net971[0:47]), .sp4_h_l_03(net1248[0:47]),
     .sp4_h_l_02(net1249[0:47]), .sp4_h_l_01(net1250[0:47]),
     .bl(bl[125:72]), .bot_op_01(bot_op_02_09[7:0]),
     .sp12_h_l_01(net1240[0:23]), .sp12_h_l_02(net1239[0:23]),
     .sp12_h_l_03(net1238[0:23]), .sp12_h_l_04(net1237[0:23]),
     .sp4_v_b_04(net1243[0:47]), .sp4_v_b_03(net1244[0:47]),
     .sp4_v_b_02(net1245[0:47]), .bnr_op_01(bnr_op_02_09[7:0]),
     .sp4_h_l_05(net1271[0:47]), .sp4_h_l_06(net1270[0:47]),
     .sp4_h_l_07(net1269[0:47]), .sp4_h_l_08(net1268[0:47]),
     .sp4_h_r_08(net989[0:47]), .sp4_h_r_07(net990[0:47]),
     .sp4_h_r_06(net991[0:47]), .sp4_h_r_05(net992[0:47]),
     .slf_op_05(net1279[0:7]), .slf_op_06(net1278[0:7]),
     .slf_op_07(net1277[0:7]), .slf_op_08(net1427[0:7]),
     .rgt_op_08(net1426[0:7]), .rgt_op_07(net998[0:7]),
     .rgt_op_06(net999[0:7]), .rgt_op_05(net1000[0:7]),
     .lft_op_08(net695[0:7]), .lft_op_07(net691[0:7]),
     .lft_op_06(net687[0:7]), .lft_op_05(net683[0:7]),
     .sp12_h_l_08(net1290[0:23]), .sp12_h_l_07(net1289[0:23]),
     .sp12_h_l_06(net1288[0:23]), .sp12_h_r_05(net1008[0:23]),
     .sp12_h_r_06(net1009[0:23]), .sp12_h_r_07(net1010[0:23]),
     .sp12_h_r_08(net1011[0:23]), .sp12_h_l_05(net1287[0:23]),
     .sp4_r_v_b_05(net1013[0:47]), .sp4_r_v_b_06(net1014[0:47]),
     .sp4_r_v_b_07(net1015[0:47]), .sp4_r_v_b_08(net1016[0:47]),
     .sp4_v_b_08(net1295[0:47]), .sp4_v_b_07(net1294[0:47]),
     .sp4_v_b_06(net1293[0:47]), .sp4_v_b_05(net1292[0:47]));
ice1f_array_LT_top I_lt_col_t06 ( .glb_netwk_to(net1021[0:7]),
     .glb_netwk_bo(net1022[0:7]), .vdd_cntl(vdd_cntl_l[127:0]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .top_op_08({slf_op_06_17[3], slf_op_06_17[2], slf_op_06_17[1],
     slf_op_06_17[0], slf_op_06_17[3], slf_op_06_17[2],
     slf_op_06_17[1], slf_op_06_17[0]}), .tnl_op_08({slf_op_05_17[3],
     slf_op_05_17[2], slf_op_05_17[1], slf_op_05_17[0],
     slf_op_05_17[3], slf_op_05_17[2], slf_op_05_17[1],
     slf_op_05_17[0]}), .tnr_op_08({tnr_op_06_16[3], tnr_op_06_16[2],
     tnr_op_06_16[1], tnr_op_06_16[0], tnr_op_06_16[3],
     tnr_op_06_16[2], tnr_op_06_16[1], tnr_op_06_16[0]}),
     .sp12_v_t_08(net1029[0:23]), .sp4_v_t_08(net1030[0:47]),
     .wl(wl_l[127:0]), .rgt_op_03(rgt_op_06_11[7:0]),
     .slf_op_02(slf_op_06_10[7:0]), .rgt_op_02(rgt_op_06_10[7:0]),
     .rgt_op_01(rgt_op_06_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net1135[0:7]), .lft_op_03(net1125[0:7]),
     .lft_op_02(net1127[0:7]), .lft_op_01(slf_op_05_09[7:0]),
     .rgt_op_04(rgt_op_06_12[7:0]), .carry_in(carry_in_06_09),
     .bnl_op_01(bnl_op_06_09[7:0]), .slf_op_04(slf_op_06_12[7:0]),
     .slf_op_03(slf_op_06_11[7:0]), .slf_op_01(slf_op_06_09[7:0]),
     .sp4_h_l_04(net1340[0:47]), .carry_out(net1420),
     .sp12_v_b__01(sp12_v_b_06_09[23:0]),
     .sp12_h_r_04(sp12_h_r_06_12[23:0]),
     .sp12_h_r_03(sp12_h_r_06_11[23:0]),
     .sp12_h_r_02(sp12_h_r_06_10[23:0]),
     .sp12_h_r_01(sp12_h_r_06_09[23:0]),
     .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_06_09[47:0]),
     .sp4_r_v_b_04(sp4_r_v_b_06_12[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_06_11[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_06_10[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_06_09[47:0]),
     .sp4_h_r_04(sp4_h_r_06_12[47:0]),
     .sp4_h_r_03(sp4_h_r_06_11[47:0]),
     .sp4_h_r_02(sp4_h_r_06_10[47:0]),
     .sp4_h_r_01(sp4_h_r_06_09[47:0]), .sp4_h_l_03(net1341[0:47]),
     .sp4_h_l_02(net1342[0:47]), .sp4_h_l_01(net1343[0:47]),
     .bl(bl[329:276]), .bot_op_01(bot_op_06_09[7:0]),
     .sp12_h_l_01(net1333[0:23]), .sp12_h_l_02(net1332[0:23]),
     .sp12_h_l_03(net1331[0:23]), .sp12_h_l_04(net1330[0:23]),
     .sp4_v_b_04(net1336[0:47]), .sp4_v_b_03(net1337[0:47]),
     .sp4_v_b_02(net1338[0:47]), .bnr_op_01(bnr_op_06_09[7:0]),
     .sp4_h_l_05(net1364[0:47]), .sp4_h_l_06(net1363[0:47]),
     .sp4_h_l_07(net1362[0:47]), .sp4_h_l_08(net1361[0:47]),
     .sp4_h_r_08(sp4_h_r_06_16[47:0]),
     .sp4_h_r_07(sp4_h_r_06_15[47:0]),
     .sp4_h_r_06(sp4_h_r_06_14[47:0]),
     .sp4_h_r_05(sp4_h_r_06_13[47:0]), .slf_op_05(slf_op_06_13[7:0]),
     .slf_op_06(slf_op_06_14[7:0]), .slf_op_07(slf_op_06_15[7:0]),
     .slf_op_08(slf_op_06_16[7:0]), .rgt_op_08(rgt_op_06_16[7:0]),
     .rgt_op_07(rgt_op_06_15[7:0]), .rgt_op_06(rgt_op_06_14[7:0]),
     .rgt_op_05(rgt_op_06_13[7:0]), .lft_op_08(net1445[0:7]),
     .lft_op_07(net1184[0:7]), .lft_op_06(net1185[0:7]),
     .lft_op_05(net1186[0:7]), .sp12_h_l_08(net1383[0:23]),
     .sp12_h_l_07(net1382[0:23]), .sp12_h_l_06(net1381[0:23]),
     .sp12_h_r_05(sp12_h_r_06_13[23:0]),
     .sp12_h_r_06(sp12_h_r_06_14[23:0]),
     .sp12_h_r_07(sp12_h_r_06_15[23:0]),
     .sp12_h_r_08(sp12_h_r_06_16[23:0]), .sp12_h_l_05(net1380[0:23]),
     .sp4_r_v_b_05(sp4_r_v_b_06_13[47:0]),
     .sp4_r_v_b_06(sp4_r_v_b_06_14[47:0]),
     .sp4_r_v_b_07(sp4_r_v_b_06_15[47:0]),
     .sp4_r_v_b_08(sp4_r_v_b_06_16[47:0]), .sp4_v_b_08(net1388[0:47]),
     .sp4_v_b_07(net1387[0:47]), .sp4_v_b_06(net1386[0:47]),
     .sp4_v_b_05(net1385[0:47]));
ice1f_array_LT_top I_lt_col_t04 ( .glb_netwk_to(net1114[0:7]),
     .glb_netwk_bo(net1405[0:7]), .vdd_cntl(vdd_cntl_l[127:0]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .top_op_08({slf_op_04_17[3], slf_op_04_17[2], slf_op_04_17[1],
     slf_op_04_17[0], slf_op_04_17[3], slf_op_04_17[2],
     slf_op_04_17[1], slf_op_04_17[0]}), .tnl_op_08({slf_op_03_17[3],
     slf_op_03_17[2], slf_op_03_17[1], slf_op_03_17[0],
     slf_op_03_17[3], slf_op_03_17[2], slf_op_03_17[1],
     slf_op_03_17[0]}), .tnr_op_08({slf_op_05_17[3], slf_op_05_17[2],
     slf_op_05_17[1], slf_op_05_17[0], slf_op_05_17[3],
     slf_op_05_17[2], slf_op_05_17[1], slf_op_05_17[0]}),
     .sp12_v_t_08(net1122[0:23]), .sp4_v_t_08(net1123[0:47]),
     .wl(wl_l[127:0]), .rgt_op_03(net1125[0:7]),
     .slf_op_02(net898[0:7]), .rgt_op_02(net1127[0:7]),
     .rgt_op_01(slf_op_05_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net949[0:7]), .lft_op_03(net939[0:7]),
     .lft_op_02(net941[0:7]), .lft_op_01(slf_op_03_09[7:0]),
     .rgt_op_04(net1135[0:7]), .carry_in(carry_in_04_09),
     .bnl_op_01(bnl_op_04_09[7:0]), .slf_op_04(net900[0:7]),
     .slf_op_03(net897[0:7]), .slf_op_01(slf_op_04_09[7:0]),
     .sp4_h_l_04(net909[0:47]), .carry_out(net1429),
     .sp12_v_b__01(sp12_v_b_04_09[23:0]), .sp12_h_r_04(net1144[0:23]),
     .sp12_h_r_03(net1145[0:23]), .sp12_h_r_02(net1146[0:23]),
     .sp12_h_r_01(net1147[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_04_09[47:0]), .sp4_r_v_b_04(net1150[0:47]),
     .sp4_r_v_b_03(net1151[0:47]), .sp4_r_v_b_02(net1152[0:47]),
     .sp4_r_v_b_01(sp4_v_b_05_09[47:0]), .sp4_h_r_04(net1154[0:47]),
     .sp4_h_r_03(net1155[0:47]), .sp4_h_r_02(net1156[0:47]),
     .sp4_h_r_01(net1157[0:47]), .sp4_h_l_03(net910[0:47]),
     .sp4_h_l_02(net911[0:47]), .sp4_h_l_01(net912[0:47]),
     .bl(bl[221:168]), .bot_op_01(bot_op_04_09[7:0]),
     .sp12_h_l_01(net883[0:23]), .sp12_h_l_02(net885[0:23]),
     .sp12_h_l_03(net844[0:23]), .sp12_h_l_04(net887[0:23]),
     .sp4_v_b_04(net860[0:47]), .sp4_v_b_03(net858[0:47]),
     .sp4_v_b_02(net856[0:47]), .bnr_op_01(bnr_op_04_09[7:0]),
     .sp4_h_l_05(net919[0:47]), .sp4_h_l_06(net917[0:47]),
     .sp4_h_l_07(net878[0:47]), .sp4_h_l_08(net879[0:47]),
     .sp4_h_r_08(net1175[0:47]), .sp4_h_r_07(net1176[0:47]),
     .sp4_h_r_06(net1177[0:47]), .sp4_h_r_05(net1178[0:47]),
     .slf_op_05(net906[0:7]), .slf_op_06(net907[0:7]),
     .slf_op_07(net894[0:7]), .slf_op_08(net895[0:7]),
     .rgt_op_08(net1445[0:7]), .rgt_op_07(net1184[0:7]),
     .rgt_op_06(net1185[0:7]), .rgt_op_05(net1186[0:7]),
     .lft_op_08(net1426[0:7]), .lft_op_07(net998[0:7]),
     .lft_op_06(net999[0:7]), .lft_op_05(net1000[0:7]),
     .sp12_h_l_08(net843[0:23]), .sp12_h_l_07(net847[0:23]),
     .sp12_h_l_06(net840[0:23]), .sp12_h_r_05(net1194[0:23]),
     .sp12_h_r_06(net1195[0:23]), .sp12_h_r_07(net1196[0:23]),
     .sp12_h_r_08(net1197[0:23]), .sp12_h_l_05(net842[0:23]),
     .sp4_r_v_b_05(net1199[0:47]), .sp4_r_v_b_06(net1200[0:47]),
     .sp4_r_v_b_07(net1201[0:47]), .sp4_r_v_b_08(net1202[0:47]),
     .sp4_v_b_08(net881[0:47]), .sp4_v_b_07(net880[0:47]),
     .sp4_v_b_06(net861[0:47]), .sp4_v_b_05(net863[0:47]));
ice1f_array_LT_top I_lt_col_t01 ( .glb_netwk_to(net1207[0:7]),
     .glb_netwk_bo(net1406[0:7]), .vdd_cntl(vdd_cntl_l[127:0]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .top_op_08({slf_op_01_17[3], slf_op_01_17[2], slf_op_01_17[1],
     slf_op_01_17[0], slf_op_01_17[3], slf_op_01_17[2],
     slf_op_01_17[1], slf_op_01_17[0]}), .tnl_op_08({tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .tnr_op_08({slf_op_02_17[3], slf_op_02_17[2], slf_op_02_17[1],
     slf_op_02_17[0], slf_op_02_17[3], slf_op_02_17[2],
     slf_op_02_17[1], slf_op_02_17[0]}), .sp12_v_t_08(net1215[0:23]),
     .sp4_v_t_08(net1216[0:47]), .wl(wl_l[127:0]),
     .rgt_op_03(net1218[0:7]), .slf_op_02(net671[0:7]),
     .rgt_op_02(net1220[0:7]), .rgt_op_01(slf_op_02_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04({slf_op_00_12[3],
     slf_op_00_12[2], slf_op_00_12[1], slf_op_00_12[0],
     slf_op_00_12[3], slf_op_00_12[2], slf_op_00_12[1],
     slf_op_00_12[0]}), .lft_op_03({slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0], slf_op_00_11[3],
     slf_op_00_11[2], slf_op_00_11[1], slf_op_00_11[0]}),
     .lft_op_02({slf_op_00_10[3], slf_op_00_10[2], slf_op_00_10[1],
     slf_op_00_10[0], slf_op_00_10[3], slf_op_00_10[2],
     slf_op_00_10[1], slf_op_00_10[0]}), .lft_op_01({slf_op_00_09[3],
     slf_op_00_09[2], slf_op_00_09[1], slf_op_00_09[0],
     slf_op_00_09[3], slf_op_00_09[2], slf_op_00_09[1],
     slf_op_00_09[0]}), .rgt_op_04(net1228[0:7]),
     .carry_in(carry_in_01_09), .bnl_op_01(bnl_op_01_09[7:0]),
     .slf_op_04(net679[0:7]), .slf_op_03(net675[0:7]),
     .slf_op_01(slf_op_01_09[7:0]), .sp4_h_l_04(net676[0:47]),
     .carry_out(net1421), .sp12_v_b__01(sp12_v_b_01_09[23:0]),
     .sp12_h_r_04(net1237[0:23]), .sp12_h_r_03(net1238[0:23]),
     .sp12_h_r_02(net1239[0:23]), .sp12_h_r_01(net1240[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_01_09[47:0]), .sp4_r_v_b_04(net1243[0:47]),
     .sp4_r_v_b_03(net1244[0:47]), .sp4_r_v_b_02(net1245[0:47]),
     .sp4_r_v_b_01(sp4_v_b_02_09[47:0]), .sp4_h_r_04(net1247[0:47]),
     .sp4_h_r_03(net1248[0:47]), .sp4_h_r_02(net1249[0:47]),
     .sp4_h_r_01(net1250[0:47]), .sp4_h_l_03(net672[0:47]),
     .sp4_h_l_02(net668[0:47]), .sp4_h_l_01(net664[0:47]),
     .bl(bl[71:18]), .bot_op_01(bot_op_01_09[7:0]),
     .sp12_h_l_01(net665[0:23]), .sp12_h_l_02(net669[0:23]),
     .sp12_h_l_03(net673[0:23]), .sp12_h_l_04(net677[0:23]),
     .sp4_v_b_04(net1460[0:47]), .sp4_v_b_03(net1475[0:47]),
     .sp4_v_b_02(net1412[0:47]), .bnr_op_01(bnr_op_01_09[7:0]),
     .sp4_h_l_05(net680[0:47]), .sp4_h_l_06(net684[0:47]),
     .sp4_h_l_07(net688[0:47]), .sp4_h_l_08(net692[0:47]),
     .sp4_h_r_08(net1268[0:47]), .sp4_h_r_07(net1269[0:47]),
     .sp4_h_r_06(net1270[0:47]), .sp4_h_r_05(net1271[0:47]),
     .slf_op_05(net683[0:7]), .slf_op_06(net687[0:7]),
     .slf_op_07(net691[0:7]), .slf_op_08(net695[0:7]),
     .rgt_op_08(net1427[0:7]), .rgt_op_07(net1277[0:7]),
     .rgt_op_06(net1278[0:7]), .rgt_op_05(net1279[0:7]),
     .lft_op_08({slf_op_00_16[3], slf_op_00_16[2], slf_op_00_16[1],
     slf_op_00_16[0], slf_op_00_16[3], slf_op_00_16[2],
     slf_op_00_16[1], slf_op_00_16[0]}), .lft_op_07({slf_op_00_15[3],
     slf_op_00_15[2], slf_op_00_15[1], slf_op_00_15[0],
     slf_op_00_15[3], slf_op_00_15[2], slf_op_00_15[1],
     slf_op_00_15[0]}), .lft_op_06({slf_op_00_14[3], slf_op_00_14[2],
     slf_op_00_14[1], slf_op_00_14[0], slf_op_00_14[3],
     slf_op_00_14[2], slf_op_00_14[1], slf_op_00_14[0]}),
     .lft_op_05({slf_op_00_13[3], slf_op_00_13[2], slf_op_00_13[1],
     slf_op_00_13[0], slf_op_00_13[3], slf_op_00_13[2],
     slf_op_00_13[1], slf_op_00_13[0]}), .sp12_h_l_08(net1424[0:23]),
     .sp12_h_l_07(net1444[0:23]), .sp12_h_l_06(net685[0:23]),
     .sp12_h_r_05(net1287[0:23]), .sp12_h_r_06(net1288[0:23]),
     .sp12_h_r_07(net1289[0:23]), .sp12_h_r_08(net1290[0:23]),
     .sp12_h_l_05(net681[0:23]), .sp4_r_v_b_05(net1292[0:47]),
     .sp4_r_v_b_06(net1293[0:47]), .sp4_r_v_b_07(net1294[0:47]),
     .sp4_r_v_b_08(net1295[0:47]), .sp4_v_b_08(net1435[0:47]),
     .sp4_v_b_07(net1441[0:47]), .sp4_v_b_06(net1413[0:47]),
     .sp4_v_b_05(net1419[0:47]));
ice1f_array_LT_top I_lt_col_t05 ( .glb_netwk_to(net1300[0:7]),
     .glb_netwk_bo(net1414[0:7]), .vdd_cntl(vdd_cntl_l[127:0]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .top_op_08({slf_op_05_17[3], slf_op_05_17[2], slf_op_05_17[1],
     slf_op_05_17[0], slf_op_05_17[3], slf_op_05_17[2],
     slf_op_05_17[1], slf_op_05_17[0]}), .tnl_op_08({slf_op_04_17[3],
     slf_op_04_17[2], slf_op_04_17[1], slf_op_04_17[0],
     slf_op_04_17[3], slf_op_04_17[2], slf_op_04_17[1],
     slf_op_04_17[0]}), .tnr_op_08({slf_op_06_17[3], slf_op_06_17[2],
     slf_op_06_17[1], slf_op_06_17[0], slf_op_06_17[3],
     slf_op_06_17[2], slf_op_06_17[1], slf_op_06_17[0]}),
     .sp12_v_t_08(net1308[0:23]), .sp4_v_t_08(net1309[0:47]),
     .wl(wl_l[127:0]), .rgt_op_03(slf_op_06_11[7:0]),
     .slf_op_02(net1127[0:7]), .rgt_op_02(slf_op_06_10[7:0]),
     .rgt_op_01(slf_op_06_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net900[0:7]), .lft_op_03(net897[0:7]),
     .lft_op_02(net898[0:7]), .lft_op_01(slf_op_04_09[7:0]),
     .rgt_op_04(slf_op_06_12[7:0]), .carry_in(carry_in_05_09),
     .bnl_op_01(bnl_op_05_09[7:0]), .slf_op_04(net1135[0:7]),
     .slf_op_03(net1125[0:7]), .slf_op_01(slf_op_05_09[7:0]),
     .sp4_h_l_04(net1154[0:47]), .carry_out(net1328),
     .sp12_v_b__01(sp12_v_b_05_09[23:0]), .sp12_h_r_04(net1330[0:23]),
     .sp12_h_r_03(net1331[0:23]), .sp12_h_r_02(net1332[0:23]),
     .sp12_h_r_01(net1333[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .sp4_v_b_01(sp4_v_b_05_09[47:0]), .sp4_r_v_b_04(net1336[0:47]),
     .sp4_r_v_b_03(net1337[0:47]), .sp4_r_v_b_02(net1338[0:47]),
     .sp4_r_v_b_01(sp4_v_b_06_09[47:0]), .sp4_h_r_04(net1340[0:47]),
     .sp4_h_r_03(net1341[0:47]), .sp4_h_r_02(net1342[0:47]),
     .sp4_h_r_01(net1343[0:47]), .sp4_h_l_03(net1155[0:47]),
     .sp4_h_l_02(net1156[0:47]), .sp4_h_l_01(net1157[0:47]),
     .bl(bl[275:222]), .bot_op_01(bot_op_05_09[7:0]),
     .sp12_h_l_01(net1147[0:23]), .sp12_h_l_02(net1146[0:23]),
     .sp12_h_l_03(net1145[0:23]), .sp12_h_l_04(net1144[0:23]),
     .sp4_v_b_04(net1150[0:47]), .sp4_v_b_03(net1151[0:47]),
     .sp4_v_b_02(net1152[0:47]), .bnr_op_01(bnr_op_05_09[7:0]),
     .sp4_h_l_05(net1178[0:47]), .sp4_h_l_06(net1177[0:47]),
     .sp4_h_l_07(net1176[0:47]), .sp4_h_l_08(net1175[0:47]),
     .sp4_h_r_08(net1361[0:47]), .sp4_h_r_07(net1362[0:47]),
     .sp4_h_r_06(net1363[0:47]), .sp4_h_r_05(net1364[0:47]),
     .slf_op_05(net1186[0:7]), .slf_op_06(net1185[0:7]),
     .slf_op_07(net1184[0:7]), .slf_op_08(net1445[0:7]),
     .rgt_op_08(slf_op_06_16[7:0]), .rgt_op_07(slf_op_06_15[7:0]),
     .rgt_op_06(slf_op_06_14[7:0]), .rgt_op_05(slf_op_06_13[7:0]),
     .lft_op_08(net895[0:7]), .lft_op_07(net894[0:7]),
     .lft_op_06(net907[0:7]), .lft_op_05(net906[0:7]),
     .sp12_h_l_08(net1197[0:23]), .sp12_h_l_07(net1196[0:23]),
     .sp12_h_l_06(net1195[0:23]), .sp12_h_r_05(net1380[0:23]),
     .sp12_h_r_06(net1381[0:23]), .sp12_h_r_07(net1382[0:23]),
     .sp12_h_r_08(net1383[0:23]), .sp12_h_l_05(net1194[0:23]),
     .sp4_r_v_b_05(net1385[0:47]), .sp4_r_v_b_06(net1386[0:47]),
     .sp4_r_v_b_07(net1387[0:47]), .sp4_r_v_b_08(net1388[0:47]),
     .sp4_v_b_08(net1202[0:47]), .sp4_v_b_07(net1201[0:47]),
     .sp4_v_b_06(net1200[0:47]), .sp4_v_b_05(net1199[0:47]));
fabric_outbuf12p I_fbuf_f0617 ( .fabric_out(net_fabric_out_06_17),
     .cout(fabric_out_06_17));
fabric_outbuf12p I_fbuf_f0009 ( .fabric_out(net_fabric_out_00_09),
     .cout(fabric_out_00_09));
fabric_outbuf12p I_fbuf_p0009 ( .fabric_out(padinlat_l_t[0]),
     .cout(padin_00_09a));
fabric_outbuf12p I_fbuf_p0617b ( .fabric_out(padinlat_t_l[11]),
     .cout(padin_06_17b));
clk_quad_buf12px8 I_clk_quadbuf_ice1fx8 ( .clko(clk_tree_drv[7:0]),
     .clki(glb_in[7:0]));

endmodule
// Library - leafcell, Cell - clk_mux2to1ice12p, View - schematic
// LAST TIME SAVED: Mar 17 10:48:45 2009
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module clk_mux2to1ice12p ( clk, cbit, cbitb, min, prog );
output  clk;

input  cbit, cbitb, prog;

input [1:0]  min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate I290 ( .in(min[0]), .out(st2), .pp(cbit), .nn(cbitb));
txgate I295 ( .in(min[1]), .out(st2), .pp(cbitb), .nn(cbit));
inv_hvt I292 ( .A(prog), .Y(progb));
inv_hvt I294 ( .A(net86), .Y(clk));
nand2_hvt I293 ( .B(progb), .A(st2), .Y(net86));

endmodule
// Library - leafcell, Cell - ice12p_clk_mux2to1, View - schematic
// LAST TIME SAVED: Jan 21 14:06:33 2009
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module ice12p_clk_mux2to1 ( gnet, bl, min0, min1, min2, min3, pgate_l,
     pgate_r, prog, reset_l, reset_r, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r );


input  prog;

output [3:0]  gnet;

inout [3:0]  bl;

input [1:0]  wl_l;
input [1:0]  pgate_r;
input [1:0]  reset_r;
input [1:0]  vdd_cntl_r;
input [1:0]  pgate_l;
input [1:0]  wl_r;
input [1:0]  vdd_cntl_l;
input [1:0]  min0;
input [1:0]  min1;
input [1:0]  reset_l;
input [1:0]  min2;
input [1:0]  min3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [7:0]  cbitb;

wire  [0:1]  l_vdd;

wire  [7:0]  cbit;



clk_mux2to1ice12p I_ckmux3 ( .prog(prog), .cbit(cbit[3]),
     .cbitb(cbitb[3]), .min(min3[1:0]), .clk(gnet[3]));
clk_mux2to1ice12p I_ckmux1 ( .prog(prog), .cbit(cbit[1]),
     .cbitb(cbitb[1]), .min(min1[1:0]), .clk(gnet[1]));
clk_mux2to1ice12p I_ckmux2 ( .prog(prog), .cbit(cbit[2]),
     .cbitb(cbitb[2]), .min(min2[1:0]), .clk(gnet[2]));
clk_mux2to1ice12p I_ckmux0 ( .prog(prog), .cbit(cbit[0]),
     .cbitb(cbitb[0]), .min(min0[1:0]), .clk(gnet[0]));
pch_hvt  vdd_cntrl_1_ ( .D(l_vdd[0]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(l_vdd[1]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl_r[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl_r[0]), .S(vdd_));
cram2x2 I_mem30 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset_l[1:0]),
     .q(cbit[3:0]), .wl(wl_l[1:0]), .r_vdd(l_vdd[0:1]),
     .pgate(pgate_l[1:0]));
cram2x2 I_mem74 ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset_r[1:0]),
     .q(cbit[7:4]), .wl(wl_r[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate_r[1:0]));

endmodule
// Library - leafcell, Cell - bram_bufferx16_2inv, View - schematic
// LAST TIME SAVED: Aug  4 12:31:20 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module bram_bufferx16_2inv ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(in), .Y(net6));

endmodule
// Library - leafcell, Cell - bram_bufferx2e, View - schematic
// LAST TIME SAVED: Jun 25 13:54:30 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module bram_bufferx2e ( out, en, in );
output  out;

input  en, in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net7), .Y(out));
nand2_hvt I193 ( .A(en), .Y(net7), .B(in));

endmodule
// Library - misc, Cell - ml_osc, View - schematic
// LAST TIME SAVED: Sep 30 17:24:55 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_osc ( clk_out, smc_osc_fsel, smc_oscen );
output  clk_out;

input  smc_oscen;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  sel_trim;



tielo I272 ( .tielo(net0104));
tielo I273 ( .tielo(net0188));
tiehi I275 ( .tiehi(net0205));
tiehi I219 ( .tiehi(net0106));
ml_osc_stage I254 ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_b_buf), .out(out_bot), .sel_trim(sel_trim[3:0]));
ml_osc_stage I255 ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_buf), .out(out_top), .sel_trim(sel_trim[3:0]));
ml_osc_logic Iosc_logic ( .sel_trim(sel_trim[3:0]),
     .smc_oscen(smc_oscen), .smc_osc_fsel(smc_osc_fsel[1:0]),
     .clkin(clk_out));
ml_dff I174 ( .R(oscen_b), .D(clkby2_b), .CLK(clk_dffin),
     .QN(clkby2_b), .Q(clkby2));
nor3_hvt I256 ( .B(net079), .Y(net075), .A(net079), .C(net079));
nor3_hvt I218 ( .B(net083), .Y(net079), .A(net083), .C(net083));
nor3_hvt I217 ( .B(net0106), .Y(net083), .A(net0106), .C(net0106));
nand3_hvt I224 ( .Y(net088), .B(net0106), .C(net0106), .A(net0106));
nand3_hvt I230 ( .Y(net092), .B(net088), .C(net088), .A(net088));
nand3_hvt I231 ( .Y(net096), .B(net092), .C(net092), .A(net092));
rppolywo_m  R18 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(net362), .PLUS(net356), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net356), .PLUS(pbias), .BULK(gnd_));
rppolywo_m  R7 ( .BULK(gnd_), .MINUS(net383), .PLUS(net366));
rppolywo_m  R2 ( .MINUS(net366), .PLUS(net362), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net437), .PLUS(net383), .BULK(gnd_));
nand2_hvt I175 ( .A(out_bot), .Y(clk_dffin), .B(out_top));
inv_hvt I222 ( .A(clkby2), .Y(clkby2_b_buf));
inv_hvt I220 ( .A(clkby2_b), .Y(clkby2_buf));
inv_hvt I176 ( .A(clkby2_b), .Y(clk_out));
inv_hvt I248 ( .A(net0104), .Y(net0226));
inv_hvt I198 ( .A(smc_oscen), .Y(oscen_b));
nch_hvt  M45 ( .D(gnd_), .B(gnd_), .G(net0188), .S(gnd_));
nch_hvt  MN31 ( .D(net437), .B(gnd_), .G(smc_oscen), .S(gnd_));
nch_hvt  MN44 ( .D(pbias), .B(gnd_), .G(net0104), .S(net371));
pch_hvt  MP77 ( .D(net371), .B(vdd_), .G(net0226), .S(pbias));
pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(net0205), .S(vdd_));
pch_hvt  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  MP41 ( .D(pbias), .B(vdd_), .G(smc_oscen), .S(vdd_));

endmodule
// Library - leafcell, Cell - bram_bank_logic_bot, View - schematic
// LAST TIME SAVED: Aug 31 18:48:17 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module bram_bank_logic_bot ( bm_sclkrw_o, bm_sdo_o, bm_sweb_o,
     bm_banksel_i, bm_sclk_i, bm_sclkrw_i, bm_sdo_i, bm_sweb_i );

input  bm_sclk_i, bm_sclkrw_i, bm_sweb_i;

output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sclkrw_o;

input [1:0]  bm_banksel_i;
input [1:0]  bm_sdo_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net25;

wire  [1:0]  net26;



bram_bufferx16_2inv I51_1_ ( .in(net26[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I51_0_ ( .in(net26[0]), .out(bm_sdo_o[0]));
leafcell_ml_dff_schematic I52_1_ ( .R(net020), .D(bm_sdo_i[1]),
     .CLK(bm_sclk_i), .QN(net25[0]), .Q(net26[1]));
leafcell_ml_dff_schematic I52_0_ ( .R(net020), .D(bm_sdo_i[0]),
     .CLK(bm_sclk_i), .QN(net25[1]), .Q(net26[0]));
bram_bufferx2e I54_1_ ( .in(bm_sweb_i), .en(bm_banksel_i[1]),
     .out(bm_sweb_o[1]));
bram_bufferx2e I54_0_ ( .in(bm_sweb_i), .en(bm_banksel_i[0]),
     .out(bm_sweb_o[0]));
bram_bufferx2e I48_1_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[1]),
     .out(bm_sclkrw_o[1]));
bram_bufferx2e I48_0_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[0]),
     .out(bm_sclkrw_o[0]));
tielo I55 ( .tielo(net020));

endmodule
// Library - leafcell, Cell - bram_hbuffer_2xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:01:06 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module bram_hbuffer_2xbank ( bm_banksel_o, bm_init_o, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;
output [3:0]  bm_sdi_o;
output [3:0]  bm_sdo_o;
output [3:0]  bm_banksel_o;

input [3:0]  bm_sdi_i;
input [3:0]  bm_banksel_i;
input [3:0]  bm_sdo_i;
input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx16_2inv I6_3_ ( .in(bm_sdi_i[3]), .out(bm_sdi_o[3]));
bram_bufferx16_2inv I6_2_ ( .in(bm_sdi_i[2]), .out(bm_sdi_o[2]));
bram_bufferx16_2inv I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx16_2inv I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx16_2inv I5 ( .in(bm_wdummymux_en_i),
     .out(bm_wdummymux_en_o));
bram_bufferx16_2inv I2_3_ ( .in(bm_sdo_i[3]), .out(bm_sdo_o[3]));
bram_bufferx16_2inv I2_2_ ( .in(bm_sdo_i[2]), .out(bm_sdo_o[2]));
bram_bufferx16_2inv I2_1_ ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I2_0_ ( .in(bm_sdo_i[0]), .out(bm_sdo_o[0]));
bram_bufferx16_2inv I13_3_ ( .in(bm_banksel_i[3]),
     .out(bm_banksel_o[3]));
bram_bufferx16_2inv I13_2_ ( .in(bm_banksel_i[2]),
     .out(bm_banksel_o[2]));
bram_bufferx16_2inv I13_1_ ( .in(bm_banksel_i[1]),
     .out(bm_banksel_o[1]));
bram_bufferx16_2inv I13_0_ ( .in(bm_banksel_i[0]),
     .out(bm_banksel_o[0]));
bram_bufferx16_2inv I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx16_2inv I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx16_2inv I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx16_2inv I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx16_2inv I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx16_2inv I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx16_2inv I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx16_2inv I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx16_2inv I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx16_2inv I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx16_2inv I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx16_2inv I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx16_2inv I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx16_2inv I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - bram_icg, View - schematic
// LAST TIME SAVED: Jun 25 14:02:00 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module bram_icg ( clkout, clk, en );
output  clkout;

input  clk, en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(net027), .Y(net014), .B(c));
inv_tri_2_hvt I7 ( .Tb(cn), .T(c), .A(net027), .Y(net023));
inv_tri_2_hvt I5 ( .Tb(c), .T(cn), .A(en), .Y(net023));
inv_hvt I391 ( .A(net014), .Y(clkout));
inv_hvt I6 ( .A(net023), .Y(net027));
inv_hvt I4 ( .A(cn), .Y(c));
inv_hvt I3 ( .A(clk), .Y(cn));

endmodule
// Library - leafcell, Cell - bram_hbuffer_dff_2xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:02:56 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module bram_hbuffer_dff_2xbank ( bm_banksel_o, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclkrw_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [3:0]  bm_sdi_o;
output [3:0]  bm_banksel_o;
output [1:0]  bm_sclk_o;
output [7:0]  bm_sa_o;
output [3:0]  bm_sdo_o;

input [7:0]  bm_sa_i;
input [3:0]  bm_sdo_i;
input [3:0]  bm_banksel_i;
input [3:0]  bm_sdi_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net102;

wire  [0:3]  net103;



tielo I23 ( .tielo(net057));
bram_icg I47 ( .en(net74), .clk(bm_sclk_i), .clkout(net61));
bram_icg I19 ( .en(net72), .clk(bm_sclk_i), .clkout(net64));
bram_bufferx16_2inv I16_3_ ( .in(net103[0]), .out(bm_sdo_o[3]));
bram_bufferx16_2inv I16_2_ ( .in(net103[1]), .out(bm_sdo_o[2]));
bram_bufferx16_2inv I16_1_ ( .in(net103[2]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I16_0_ ( .in(net103[3]), .out(bm_sdo_o[0]));
bram_bufferx4 I6_3_ ( .in(bm_sdi_i[3]), .out(bm_sdi_o[3]));
bram_bufferx4 I6_2_ ( .in(bm_sdi_i[2]), .out(bm_sdi_o[2]));
bram_bufferx4 I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx4 I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx4 I22 ( .in(net64), .out(bm_sclk_o[1]));
bram_bufferx4 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx4 I13_3_ ( .in(bm_banksel_i[3]), .out(bm_banksel_o[3]));
bram_bufferx4 I13_2_ ( .in(bm_banksel_i[2]), .out(bm_banksel_o[2]));
bram_bufferx4 I13_1_ ( .in(bm_banksel_i[1]), .out(bm_banksel_o[1]));
bram_bufferx4 I13_0_ ( .in(bm_banksel_i[0]), .out(bm_banksel_o[0]));
bram_bufferx4 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx4 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx4 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx4 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx4 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx4 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx4 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx4 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx4 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx4 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx4 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx4 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx4 I18 ( .in(net61), .out(bm_sclk_o[0]));
bram_bufferx4 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));
leafcell_ml_dff_schematic I48_3_ ( .R(net057), .D(bm_sdo_i[3]),
     .CLK(bm_sclk_i), .QN(net102[0]), .Q(net103[0]));
leafcell_ml_dff_schematic I48_2_ ( .R(net057), .D(bm_sdo_i[2]),
     .CLK(bm_sclk_i), .QN(net102[1]), .Q(net103[1]));
leafcell_ml_dff_schematic I48_1_ ( .R(net057), .D(bm_sdo_i[1]),
     .CLK(bm_sclk_i), .QN(net102[2]), .Q(net103[2]));
leafcell_ml_dff_schematic I48_0_ ( .R(net057), .D(bm_sdo_i[0]),
     .CLK(bm_sclk_i), .QN(net102[3]), .Q(net103[3]));
nor2_hvt I20 ( .A(bm_banksel_i[2]), .B(bm_banksel_i[3]), .Y(net67));
nor2_hvt I49 ( .A(bm_banksel_i[0]), .B(bm_banksel_i[1]), .Y(net70));
inv_hvt I21 ( .A(net67), .Y(net72));
inv_hvt I17 ( .A(net70), .Y(net74));

endmodule
// Library - leafcell, Cell - bram_hbuffer_1xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:50:36 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module bram_hbuffer_1xbank ( bm_banksel_o, bm_init_o, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;
output [1:0]  bm_sdi_o;
output [1:0]  bm_banksel_o;
output [1:0]  bm_sdo_o;

input [1:0]  bm_sdo_i;
input [1:0]  bm_banksel_i;
input [1:0]  bm_sdi_i;
input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx16_2inv I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx16_2inv I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx16_2inv I5 ( .in(bm_wdummymux_en_i),
     .out(bm_wdummymux_en_o));
bram_bufferx16_2inv I2_1_ ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I2_0_ ( .in(bm_sdo_i[0]), .out(bm_sdo_o[0]));
bram_bufferx16_2inv I13_1_ ( .in(bm_banksel_i[1]),
     .out(bm_banksel_o[1]));
bram_bufferx16_2inv I13_0_ ( .in(bm_banksel_i[0]),
     .out(bm_banksel_o[0]));
bram_bufferx16_2inv I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx16_2inv I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx16_2inv I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx16_2inv I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx16_2inv I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx16_2inv I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx16_2inv I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx16_2inv I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx16_2inv I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx16_2inv I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx16_2inv I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx16_2inv I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx16_2inv I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx16_2inv I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - ice1f_quad_x4, View - schematic
// LAST TIME SAVED: Aug 15 14:59:41 2009
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module ice1f_quad_x4 ( bm_sdo_o, cf_b, cf_l, cf_r, cf_t,
     fabric_out_12_00_wb, fabric_out_13_01_wb_sel0,
     fabric_out_13_02_wb_sel1, padeb_b, padeb_l, padeb_r, padeb_t,
     pado_b, pado_l, pado_r, pado_t, sdo_pad, spi_ss_in_b, spi_ss_in_l,
     spi_ss_in_r, bl_bot, bl_top, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en, ceb,
     end_of_startup_b, end_of_startup_l, end_of_startup_r,
     end_of_startup_t, hiz_b, last_rsr, mode, padin_b, padin_l,
     padin_r, padin_t, pgate_l, pgate_r, prog, purst, r, reset_b_l,
     reset_b_r, sdi_pad, shift, spioeb_b, spioeb_l, spiout_b, spiout_l,
     spiout_r, tclk, tiegnd, tievdd, update, vdd_cntl_l, vdd_cntl_r,
     wl_l, wl_r );
output  fabric_out_12_00_wb, fabric_out_13_01_wb_sel0,
     fabric_out_13_02_wb_sel1, sdo_pad;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en, ceb, hiz_b, last_rsr, mode,
     prog, purst, r, sdi_pad, shift, tclk, tiegnd, tievdd, update;

output [15:0]  spi_ss_in_l;
output [3:0]  bm_sdo_o;
output [23:12]  spi_ss_in_b;
output [31:0]  spi_ss_in_r;
output [23:0]  padeb_b;
output [287:0]  cf_b;
output [23:0]  padeb_t;
output [383:0]  cf_l;
output [23:0]  pado_b;
output [23:0]  pado_t;
output [20:0]  padeb_r;
output [20:0]  pado_r;
output [25:0]  padeb_l;
output [383:0]  cf_r;
output [25:0]  pado_l;
output [287:0]  cf_t;

inout [663:0]  bl_bot;
inout [663:0]  bl_top;

input [23:12]  spiout_b;
input [3:0]  bm_banksel_i;
input [15:0]  spiout_r;
input [3:0]  bm_sdi_i;
input [15:0]  spioeb_l;
input [15:0]  spiout_l;
input [287:0]  wl_r;
input [23:12]  spioeb_b;
input [287:0]  wl_l;
input [23:0]  padin_b;
input [16:1]  end_of_startup_l;
input [12:7]  end_of_startup_b;
input [7:0]  bm_sa_i;
input [287:0]  vdd_cntl_r;
input [12:1]  end_of_startup_t;
input [25:0]  padin_l;
input [287:0]  pgate_r;
input [16:1]  end_of_startup_r;
input [287:0]  reset_b_r;
input [20:0]  padin_r;
input [287:0]  vdd_cntl_l;
input [287:0]  pgate_l;
input [287:0]  reset_b_l;
input [23:0]  padin_t;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  slf_op_11_08;

wire  [7:0]  slf_op_06_14;

wire  [0:23]  net729;

wire  [0:23]  net595;

wire  [0:23]  net1031;

wire  [0:23]  net628;

wire  [0:23]  net1030;

wire  [0:1]  net835;

wire  [0:23]  net735;

wire  [0:23]  net592;

wire  [0:47]  net556;

wire  [0:7]  net689;

wire  [0:1]  net1273;

wire  [0:23]  net596;

wire  [0:1]  net664;

wire  [0:23]  net590;

wire  [7:0]  slf_op_10_08;

wire  [7:0]  slf_op_06_02;

wire  [0:23]  net597;

wire  [3:0]  slf_op_07_17;

wire  [0:3]  net1250;

wire  [0:47]  net727;

wire  [0:47]  net739;

wire  [0:47]  net558;

wire  [0:15]  net598;

wire  [0:7]  net1008;

wire  [0:15]  net555;

wire  [0:47]  net1076;

wire  [7:0]  slf_op_04_08;

wire  [7:0]  slf_op_07_07;

wire  [0:23]  net1081;

wire  [0:47]  net612;

wire  [7:0]  slf_op_07_01;

wire  [0:23]  net753;

wire  [7:0]  slf_op_04_09;

wire  [0:7]  net856;

wire  [7:0]  slf_op_06_11;

wire  [0:7]  net1257;

wire  [0:47]  net587;

wire  [7:0]  slf_op_07_06;

wire  [0:47]  net751;

wire  [7:0]  slf_op_06_09;

wire  [0:47]  net1079;

wire  [7:0]  slf_op_06_07;

wire  [0:7]  net1279;

wire  [0:47]  net588;

wire  [0:15]  net1055;

wire  [0:23]  net1028;

wire  [1:0]  bm_bank10_banksel_o;

wire  [3:0]  slf_op_13_08;

wire  [0:47]  net1090;

wire  [0:23]  net627;

wire  [0:23]  net625;

wire  [7:0]  slf_op_12_08;

wire  [0:47]  net613;

wire  [0:3]  net1245;

wire  [7:0]  slf_op_06_08;

wire  [7:0]  slf_op_07_02;

wire  [0:23]  net593;

wire  [0:23]  net1033;

wire  [0:23]  net626;

wire  [0:47]  net583;

wire  [7:0]  slf_op_07_08;

wire  [0:23]  net624;

wire  [0:47]  net550;

wire  [7:0]  slf_op_07_09;

wire  [0:47]  net616;

wire  [7:0]  slf_op_08_09;

wire  [0:47]  net1068;

wire  [1:0]  bm_sclkrw_b2_o;

wire  [0:47]  net1077;

wire  [7:0]  slf_op_03_08;

wire  [7:0]  slf_op_06_15;

wire  [0:3]  net1246;

wire  [0:23]  net1034;

wire  [0:47]  net611;

wire  [0:23]  net594;

wire  [0:23]  net747;

wire  [0:47]  net1075;

wire  [7:0]  gclk;

wire  [3:0]  slf_op_06_17;

wire  [0:1]  net685;

wire  [7:0]  slf_op_01_08;

wire  [0:1]  net667;

wire  [0:47]  net561;

wire  [7:0]  slf_op_05_08;

wire  [7:0]  slf_op_01_09;

wire  [0:23]  net758;

wire  [0:47]  net549;

wire  [3:0]  slf_op_00_09;

wire  [7:0]  slf_op_10_09;

wire  [0:47]  net615;

wire  [0:47]  net589;

wire  [3:0]  slf_op_13_09;

wire  [0:47]  net1091;

wire  [0:1]  net852;

wire  [0:47]  net1080;

wire  [0:47]  net585;

wire  [0:23]  net552;

wire  [7:0]  slf_op_07_11;

wire  [0:47]  net1089;

wire  [7:0]  slf_op_06_16;

wire  [7:0]  slf_op_09_08;

wire  [0:47]  net584;

wire  [1:0]  bm_sdi_b0_o;

wire  [0:1]  net1204;

wire  [3:0]  bm_bank30_sdo_i;

wire  [7:0]  slf_op_07_12;

wire  [0:1]  net1272;

wire  [0:47]  net1112;

wire  [0:23]  net1029;

wire  [7:0]  slf_op_12_09;

wire  [7:0]  slf_op_06_13;

wire  [0:1]  net668;

wire  [0:47]  net756;

wire  [0:23]  net741;

wire  [0:47]  net745;

wire  [0:7]  net1233;

wire  [0:47]  net586;

wire  [0:1]  net1255;

wire  [0:47]  net1102;

wire  [0:7]  net670;

wire  [7:0]  slf_op_07_05;

wire  [0:47]  net582;

wire  [0:47]  net1094;

wire  [1:0]  bm_sdi_b2_o;

wire  [7:0]  slf_op_07_13;

wire  [7:0]  slf_op_07_14;

wire  [7:0]  bm_sa_b1_o;

wire  [7:0]  slf_op_11_09;

wire  [0:1]  net831;

wire  [0:23]  net591;

wire  [7:0]  slf_op_06_01;

wire  [0:47]  net614;

wire  [0:47]  net560;

wire  [7:0]  slf_op_06_03;

wire  [7:0]  slf_op_03_09;

wire  [7:0]  slf_op_07_04;

wire  [7:0]  slf_op_02_08;

wire  [0:15]  net701;

wire  [1:0]  bm_sclkrw_b0_o;

wire  [1:0]  bm_sweb_b2_o;

wire  [3:0]  bm_bank30_sdi_o;

wire  [0:47]  net559;

wire  [0:47]  net557;

wire  [7:0]  slf_op_02_09;

wire  [3:0]  slf_op_06_00;

wire  [7:0]  slf_op_06_10;

wire  [1:0]  bm_bank30_sclk_o;

wire  [3:0]  bm_bank30_banksel_o;

wire  [7:0]  slf_op_07_16;

wire  [3:0]  slf_op_07_00;

wire  [7:0]  slf_op_06_12;

wire  [0:47]  net1078;

wire  [0:23]  net1032;

wire  [7:0]  slf_op_05_09;

wire  [7:0]  slf_op_07_10;

wire  [7:0]  slf_op_07_15;

wire  [0:47]  net733;

wire  [0:47]  net1092;

wire  [0:47]  net1093;

wire  [7:0]  slf_op_09_09;

wire  [7:0]  slf_op_08_08;

wire  [7:0]  slf_op_07_03;

wire  [3:0]  slf_op_00_08;

wire  [7:0]  slf_op_06_06;

wire  [1:0]  bm_sweb_b0_o;

wire  [7:0]  slf_op_06_05;

wire  [7:0]  slf_op_06_04;



// nmoscap_25  C0 ( .MINUS(gnd_), .PLUS(vdd_));
// nmoscap_25  C1 ( .MINUS(gnd_), .PLUS(vdd_));
// nmoscap_25  C2 ( .MINUS(gnd_), .PLUS(vdd_));
// nmoscap_25  C3 ( .MINUS(gnd_), .PLUS(vdd_));
// nmoscap_25  C4 ( .MINUS(gnd_), .PLUS(vdd_));
ice1f_cram_row142col4 I_ice1f_cram_row142col4top (
     .pgate_l(pgate_l[287:146]), .reset_l(reset_b_l[287:146]),
     .vdd_cntl_l(vdd_cntl_l[287:146]), .wl_l(wl_l[287:146]),
     .pgate_r(pgate_r[287:146]), .reset_r(reset_b_r[287:146]),
     .vdd_cntl_r(vdd_cntl_r[287:146]), .wl_r(wl_r[287:146]),
     .bl(bl_top[333:330]));
ice1f_cram_row142col4 I_ice1f_cram_row142col4bot (
     .bl(bl_bot[333:330]), .pgate_l(pgate_l[141:0]),
     .reset_l(reset_b_l[141:0]), .vdd_cntl_l(vdd_cntl_l[141:0]),
     .wl_l(wl_l[141:0]), .pgate_r(pgate_r[141:0]),
     .reset_r(reset_b_r[141:0]), .vdd_cntl_r(vdd_cntl_r[141:0]),
     .wl_r(wl_r[141:0]));
ice1f_quad_bl I_quad_bl_ice1f ( .padeb_l_b(padeb_l[13:0]),
     .pado_l_b(pado_l[13:0]), .padin_l_b(padin_l[13:0]),
     .padeb_b_l(padeb_b[11:0]), .pado_b_l(pado_b[11:0]),
     .padin_b_l(padin_b[11:0]), .carry_out_01_08(carry_io_01_0809),
     .carry_out_02_08(carry_io_02_0809),
     .carry_out_04_08(carry_io_04_0809),
     .carry_out_05_08(carry_io_05_0809),
     .carry_out_06_08(carry_io_06_0809),
     .fabric_out_05_00(fabric_out_05_00_bicegate),
     .sp4_h_r_06_07(net549[0:47]), .sp4_h_r_06_08(net550[0:47]),
     .fabric_out_00_08(fabric_out_00_08),
     .sp12_v_t_05_08(net552[0:23]), .padin_00_08b(padin_0008b_ck),
     .fabric_out_00_07(fabric_out_00_07_licegate),
     .sp4_h_r_06_00(net555[0:15]), .sp4_h_r_06_06(net556[0:47]),
     .sp4_h_r_06_05(net557[0:47]), .sp4_h_r_06_04(net558[0:47]),
     .sp4_h_r_06_03(net559[0:47]), .sp4_h_r_06_02(net560[0:47]),
     .sp4_h_r_06_01(net561[0:47]), .slf_op_06_07(slf_op_06_07[7:0]),
     .slf_op_06_06(slf_op_06_06[7:0]),
     .slf_op_06_05(slf_op_06_05[7:0]),
     .slf_op_06_04(slf_op_06_04[7:0]),
     .slf_op_06_03(slf_op_06_03[7:0]),
     .slf_op_06_02(slf_op_06_02[7:0]),
     .slf_op_06_01(slf_op_06_01[7:0]),
     .slf_op_06_00(slf_op_06_00[3:0]),
     .tnr_op_06_00(slf_op_07_01[7:0]),
     .rgt_op_06_08(slf_op_07_08[7:0]),
     .rgt_op_06_07(slf_op_07_07[7:0]),
     .rgt_op_06_06(slf_op_07_06[7:0]),
     .rgt_op_06_05(slf_op_07_05[7:0]),
     .rgt_op_06_04(slf_op_07_04[7:0]),
     .rgt_op_06_03(slf_op_07_03[7:0]),
     .rgt_op_06_02(slf_op_07_02[7:0]),
     .rgt_op_06_01(slf_op_07_01[7:0]),
     .bnr_op_06_01(slf_op_07_00[3:0]),
     .fabric_out_06_00(fabric_out_06_00),
     .padin_06_00b(padin_0600b_ck), .sp4_r_v_b_06_08(net582[0:47]),
     .sp4_r_v_b_06_07(net583[0:47]), .sp4_r_v_b_06_06(net584[0:47]),
     .sp4_r_v_b_06_05(net585[0:47]), .sp4_r_v_b_06_04(net586[0:47]),
     .sp4_r_v_b_06_03(net587[0:47]), .sp4_r_v_b_06_02(net588[0:47]),
     .sp4_r_v_b_06_01(net589[0:47]), .sp12_h_r_06_08(net590[0:23]),
     .sp12_h_r_06_07(net591[0:23]), .sp12_h_r_06_06(net592[0:23]),
     .sp12_h_r_06_05(net593[0:23]), .sp12_h_r_06_04(net594[0:23]),
     .sp12_h_r_06_03(net595[0:23]), .sp12_h_r_06_02(net596[0:23]),
     .sp12_h_r_06_01(net597[0:23]), .sp4_v_t_00_08(net598[0:15]),
     .slf_op_00_08(slf_op_00_08[3:0]),
     .slf_op_01_08(slf_op_01_08[7:0]),
     .slf_op_02_08(slf_op_02_08[7:0]),
     .slf_op_03_08(slf_op_03_08[7:0]),
     .slf_op_04_08(slf_op_04_08[7:0]),
     .slf_op_05_08(slf_op_05_08[7:0]), .tnl_op_01_08({slf_op_00_09[3],
     slf_op_00_09[2], slf_op_00_09[1], slf_op_00_09[0],
     slf_op_00_09[3], slf_op_00_09[2], slf_op_00_09[1],
     slf_op_00_09[0]}), .tnl_op_02_08(slf_op_01_09[7:0]),
     .tnl_op_03_08(slf_op_02_09[7:0]),
     .tnl_op_04_08(slf_op_03_09[7:0]),
     .tnl_op_05_08(slf_op_04_09[7:0]),
     .tnl_op_06_08(slf_op_05_09[7:0]), .sp4_v_t_01_08(net611[0:47]),
     .sp4_v_t_02_08(net612[0:47]), .sp4_v_t_03_08(net613[0:47]),
     .sp4_v_t_04_08(net614[0:47]), .sp4_v_t_05_08(net615[0:47]),
     .sp4_v_t_06_08(net616[0:47]), .slf_op_06_08(slf_op_06_08[7:0]),
     .top_op_01_08(slf_op_01_09[7:0]),
     .top_op_02_08(slf_op_02_09[7:0]),
     .top_op_03_08(slf_op_03_09[7:0]),
     .top_op_04_08(slf_op_04_09[7:0]),
     .top_op_05_08(slf_op_05_09[7:0]),
     .top_op_06_08(slf_op_06_09[7:0]), .sp12_v_t_01_08(net624[0:23]),
     .sp12_v_t_02_08(net625[0:23]), .sp12_v_t_03_08(net626[0:23]),
     .sp12_v_t_04_08(net627[0:23]), .sp12_v_t_06_08(net628[0:23]),
     .tnr_op_00_08(slf_op_01_09[7:0]),
     .tnr_op_01_08(slf_op_02_09[7:0]),
     .tnr_op_02_08(slf_op_03_09[7:0]),
     .tnr_op_03_08(slf_op_04_09[7:0]),
     .tnr_op_04_08(slf_op_05_09[7:0]),
     .tnr_op_05_08(slf_op_06_09[7:0]),
     .tnr_op_06_08(slf_op_07_09[7:0]), .cf_b_l(cf_b[143:0]),
     .bl(bl_bot[329:0]), .reset_b_l(reset_b_l[143:0]),
     .pgate_l(pgate_l[143:0]), .vdd_cntl_l(vdd_cntl_l[143:0]),
     .wl_l(wl_l[143:0]), .end_of_startup_lft_b(end_of_startup_l[8:1]),
     .cf_l(cf_l[191:0]), .spi_ss_in_l(spi_ss_in_l[15:0]),
     .spiout_l(spiout_l[15:0]), .spioeb_l(spioeb_l[15:0]),
     .hold_b_l(fabric_out_05_00_bicegate),
     .hold_l_b(fabric_out_00_07_licegate), .update_i(net649),
     .tievdd(tievdd), .tiegnd(tiegnd), .tclk_i(tclkio_ml),
     .shift_i(net653), .sdi(sdio_ml), .r_i(net655), .purst(purst),
     .prog(prog), .mode_i(net658), .hiz_b_i(net659),
     .glb_in(gclk[7:0]), .ceb_i(net661), .bs_en_i(net662),
     .bm_wdummymux_en_i(net663), .bm_sweb_i(net664[0:1]),
     .bm_sreb_i(net665), .bm_sdo_i({bm_sdo_b1_o, bm_sdi_b0_o[0]}),
     .bm_sdi_i(net667[0:1]), .bm_sclkrw_i(net668[0:1]),
     .bm_sclk_i(net669), .bm_sa_i(net670[0:7]),
     .bm_rcapmux_en_i(net671), .bm_init_i(net672), .update_o(net673),
     .tclk_o(tclkio_mb), .shift_o(net675), .sdo(sdio_mb), .r_o(net677),
     .mode_o(net678), .hiz_b_o(net679), .ceb_o(net680),
     .bs_en_o(net681), .bm_wdummymux_en_o(net682),
     .bm_sweb_o(bm_sweb_b0_o[1:0]), .bm_sreb_o(net684),
     .bm_sdo_o(net685[0:1]), .bm_sdi_o(bm_sdi_b0_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_b0_o[1:0]), .bm_sclk_o(net688),
     .bm_sa_o(net689[0:7]), .bm_rcapmux_en_o(net690),
     .bm_init_o(net691));
ice1f_quad_br I_quad_br_ice1f ( .padin_b_r(padin_b[23:12]),
     .pado_b_r(pado_b[23:12]), .padeb_b_r(padeb_b[23:12]),
     .padeb_r_b(padeb_r[8:0]), .pado_r_b(pado_r[8:0]),
     .padin_r_b(padin_r[8:0]), .spi_ss_in_b(spi_ss_in_b[23:12]),
     .spiout(spiout_b[23:12]), .spioeb(spioeb_b[23:12]),
     .sp4_v_t_13_08(net701[0:15]), .carry_out_07_08(carry_io_07_0809),
     .carry_out_12_08(carry_io_12_0809),
     .carry_out_11_08(carry_io_11_0809),
     .carry_out_09_08(carry_io_09_0809),
     .carry_out_08_08(carry_io_08_0809),
     .fabric_out_13_02(fabric_out_13_02_wb_sel1),
     .fabric_out_13_01(fabric_out_13_01_wb_sel0),
     .fabric_out_12_00(fabric_out_12_00_wb),
     .padin_13_08b(padin_1308b_ck),
     .fabric_out_13_08(fabric_out_13_08),
     .slf_op_13_08(slf_op_13_08[3:0]), .spi_ss_in_r(spi_ss_in_r[15:0]),
     .spiout_r(spiout_r[15:0]), .spioeb_r({tievdd, tievdd, tievdd,
     tiegnd, tievdd, tiegnd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd}),
     .pgate_r(pgate_r[143:0]), .reset_b_r(reset_b_r[143:0]),
     .wl_r(wl_r[143:0]), .vdd_cntl_r(vdd_cntl_r[143:0]),
     .cf_b(cf_b[287:144]), .bl(bl_bot[663:334]),
     .end_of_startup_bot_r(end_of_startup_b[12:7]),
     .end_of_startup_rgt_b(end_of_startup_r[8:1]), .cf_r(cf_r[191:0]),
     .tnl_op_12_08(slf_op_11_09[7:0]),
     .slf_op_12_08(slf_op_12_08[7:0]), .sp4_v_t_12_08(net727[0:47]),
     .top_op_12_08(slf_op_12_09[7:0]), .sp12_v_t_12_08(net729[0:23]),
     .tnr_op_12_08({slf_op_13_09[3], slf_op_13_09[2], slf_op_13_09[1],
     slf_op_13_09[0], slf_op_13_09[3], slf_op_13_09[2],
     slf_op_13_09[1], slf_op_13_09[0]}),
     .tnl_op_11_08(slf_op_10_09[7:0]),
     .slf_op_11_08(slf_op_11_08[7:0]), .sp4_v_t_11_08(net733[0:47]),
     .top_op_11_08(slf_op_11_09[7:0]), .sp12_v_t_11_08(net735[0:23]),
     .tnr_op_11_08(slf_op_12_09[7:0]),
     .tnl_op_10_08(slf_op_09_09[7:0]),
     .slf_op_10_08(slf_op_10_08[7:0]), .sp4_v_t_10_08(net739[0:47]),
     .top_op_10_08(slf_op_10_09[7:0]), .sp12_v_t_10_08(net741[0:23]),
     .tnr_op_10_08(slf_op_11_09[7:0]),
     .tnl_op_09_08(slf_op_08_09[7:0]),
     .slf_op_09_08(slf_op_09_08[7:0]), .sp4_v_t_09_08(net745[0:47]),
     .top_op_09_08(slf_op_09_09[7:0]), .sp12_v_t_09_08(net747[0:23]),
     .tnr_op_09_08(slf_op_10_09[7:0]),
     .tnl_op_08_08(slf_op_07_09[7:0]),
     .slf_op_08_08(slf_op_08_08[7:0]), .sp4_v_t_08_08(net751[0:47]),
     .top_op_08_08(slf_op_08_09[7:0]), .sp12_v_t_08_08(net753[0:23]),
     .tnr_op_08_08(slf_op_09_09[7:0]),
     .slf_op_07_08(slf_op_07_08[7:0]), .sp4_v_t_07_08(net756[0:47]),
     .top_op_07_08(slf_op_07_09[7:0]), .sp12_v_t_07_08(net758[0:23]),
     .tnr_op_07_08(slf_op_08_09[7:0]),
     .tnl_op_07_08(slf_op_06_09[7:0]), .sp4_h_l_07_00(net555[0:15]),
     .sp4_h_l_07_08(net550[0:47]), .sp4_h_l_07_07(net549[0:47]),
     .sp4_h_l_07_06(net556[0:47]), .sp4_h_l_07_05(net557[0:47]),
     .sp4_h_l_07_04(net558[0:47]), .sp4_h_l_07_03(net559[0:47]),
     .sp4_h_l_07_02(net560[0:47]), .sp4_h_l_07_01(net561[0:47]),
     .rgt_op_07_08(slf_op_06_08[7:0]),
     .rgt_op_07_07(slf_op_06_07[7:0]),
     .rgt_op_07_06(slf_op_06_06[7:0]),
     .rgt_op_07_05(slf_op_06_05[7:0]),
     .rgt_op_07_04(slf_op_06_04[7:0]),
     .rgt_op_07_03(slf_op_06_03[7:0]),
     .rgt_op_07_02(slf_op_06_02[7:0]),
     .rgt_op_07_01(slf_op_06_01[7:0]),
     .bnl_op_07_01(slf_op_06_00[3:0]),
     .slf_op_07_01(slf_op_07_01[7:0]),
     .slf_op_07_07(slf_op_07_07[7:0]),
     .slf_op_07_06(slf_op_07_06[7:0]),
     .slf_op_07_05(slf_op_07_05[7:0]),
     .slf_op_07_04(slf_op_07_04[7:0]),
     .slf_op_07_03(slf_op_07_03[7:0]),
     .slf_op_07_02(slf_op_07_02[7:0]),
     .slf_op_07_00(slf_op_07_00[3:0]), .sp4_v_b_07_08(net582[0:47]),
     .sp4_v_b_07_07(net583[0:47]), .sp4_v_b_07_06(net584[0:47]),
     .sp4_v_b_07_05(net585[0:47]), .sp4_v_b_07_04(net586[0:47]),
     .sp4_v_b_07_03(net587[0:47]), .sp4_v_b_07_02(net588[0:47]),
     .sp4_v_b_07_01(net589[0:47]), .fabric_out_07_00(fabric_out_07_00),
     .padin_07_00a(padin_0700a_ck), .sp12_h_l_07_08(net590[0:23]),
     .sp12_h_l_07_07(net591[0:23]), .sp12_h_l_07_06(net592[0:23]),
     .sp12_h_l_07_05(net593[0:23]), .sp12_h_l_07_04(net594[0:23]),
     .sp12_h_l_07_03(net595[0:23]), .sp12_h_l_07_02(net596[0:23]),
     .sp12_h_l_07_01(net597[0:23]), .update_mi(update), .tclk_mi(tclk),
     .shift_mi(shift), .sdi_pad(sdi_pad), .r_mi(r), .mode_mi(mode),
     .hold_r_b(fabric_out_13_10_ricegate),
     .hold_b_r(fabric_out_05_00_bicegate), .hiz_b_mi(hiz_b),
     .ceb_mi(ceb), .bs_en_mi(bs_en), .sdo_pad(sdo_pad),
     .update_i(net673), .tiegnd(tiegnd), .tclk_i(tclkio_mb),
     .shift_i(net675), .sdi(sdio_mb), .r_i(net677), .purst(purst),
     .prog(prog), .mode_i(net678), .hiz_b_i(net679),
     .glb_in(gclk[7:0]), .ceb_i(net680), .bs_en_i(net681),
     .bm_wdummymux_en_i(net1283), .bm_sweb_i(net831[0:1]),
     .bm_sreb_i(net1276), .bm_sdo_i({bm_sdo_b3_o, bm_sdi_b2_o[0]}),
     .bm_sdi_i(bm_bank30_sdi_o[3:2]), .bm_sclkrw_i(net835[0:1]),
     .bm_sclk_i(bm_bank30_sclk_o[1]), .bm_sa_i(net1279[0:7]),
     .bm_rcapmux_en_i(net1282), .bm_init_i(net1280), .update_o(net840),
     .tclk_o(tclkio_mr), .shift_o(net842), .sdo(sdio_mr), .r_o(net844),
     .mode_o(net845), .hiz_b_o(net846), .ceb_o(net847),
     .bs_en_o(net848), .bm_wdummymux_en_o(net849),
     .bm_sweb_o(bm_sweb_b2_o[1:0]), .bm_sreb_o(net851),
     .bm_sdo_o(net852[0:1]), .bm_sdi_o(bm_sdi_b2_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_b2_o[1:0]), .bm_sclk_o(net855),
     .bm_sa_o(net856[0:7]), .bm_rcapmux_en_o(net857),
     .bm_init_o(net858));
ice1f_quad_tr I_quad_tr_ice1f ( .padin_r(padin_r[20:9]),
     .pado_r(pado_r[20:9]), .padeb_r(padeb_r[20:9]),
     .padin_t_r(padin_t[23:12]), .padeb_t_r(padeb_t[23:12]),
     .pado_t_r(pado_t[23:12]),
     .fabric_out_08_17(fabric_out_08_17_ticegate),
     .fabric_out_13_09(fabric_out_13_09),
     .fabric_out_07_17(fabric_out_07_17),
     .padin_13_09a(padin_1309a_ck), .padin_07_17a(padin_0717a_ck),
     .fabric_out_13_10(fabric_out_13_10_ricegate),
     .bnl_op_07_09(slf_op_06_08[7:0]),
     .bnl_op_13_09(slf_op_12_08[7:0]),
     .slf_op_13_09(slf_op_13_09[3:0]),
     .end_of_startup_top_r(end_of_startup_t[12:7]),
     .spi_ss_in_r_t(spi_ss_in_r[31:16]), .cf_r(cf_r[383:192]),
     .end_of_startup_rgt_t(end_of_startup_r[16:9]),
     .sp4_h_l_07_17(net1055[0:15]), .slf_op_07_17(slf_op_07_17[3:0]),
     .tnl_op_07_16(slf_op_06_17[3:0]), .cf_t(cf_t[287:144]),
     .carry_in_12_09(carry_io_12_0809),
     .carry_in_11_09(carry_io_11_0809),
     .carry_in_09_09(carry_io_09_0809),
     .carry_in_08_09(carry_io_08_0809),
     .carry_in_07_09(carry_io_07_0809), .pgate_r(pgate_r[287:144]),
     .reset_b_r(reset_b_r[287:144]), .vdd_cntl_r(vdd_cntl_r[287:144]),
     .wl_r(wl_r[287:144]), .sp4_h_r_13_09(net701[0:15]),
     .bl(bl_top[663:334]), .lft_op_07_10(slf_op_06_10[7:0]),
     .slf_op_07_10(slf_op_07_10[7:0]), .sp12_h_l_07_10(net1034[0:23]),
     .sp4_v_b_07_10(net1080[0:47]), .sp4_h_l_07_10(net1094[0:47]),
     .lft_op_07_11(slf_op_06_11[7:0]),
     .slf_op_07_11(slf_op_07_11[7:0]), .sp12_h_l_07_11(net1033[0:23]),
     .sp4_v_b_07_11(net1079[0:47]), .sp4_h_l_07_11(net1093[0:47]),
     .lft_op_07_12(slf_op_06_12[7:0]),
     .slf_op_07_12(slf_op_07_12[7:0]), .sp12_h_l_07_12(net1032[0:23]),
     .sp4_v_b_07_12(net1078[0:47]), .sp4_h_l_07_12(net1092[0:47]),
     .lft_op_07_13(slf_op_06_13[7:0]),
     .slf_op_07_13(slf_op_07_13[7:0]), .sp12_h_l_07_13(net1031[0:23]),
     .sp4_v_b_07_13(net1077[0:47]), .sp4_h_l_07_13(net1091[0:47]),
     .lft_op_07_14(slf_op_06_14[7:0]),
     .slf_op_07_14(slf_op_07_14[7:0]), .sp12_h_l_07_14(net1030[0:23]),
     .sp4_v_b_07_14(net1076[0:47]), .sp4_h_l_07_14(net1090[0:47]),
     .lft_op_07_15(slf_op_06_15[7:0]),
     .slf_op_07_15(slf_op_07_15[7:0]), .sp12_h_l_07_15(net1029[0:23]),
     .sp4_v_b_07_15(net1075[0:47]), .sp4_h_l_07_15(net1089[0:47]),
     .lft_op_07_16(slf_op_06_16[7:0]),
     .slf_op_07_16(slf_op_07_16[7:0]), .sp12_h_l_07_16(net1028[0:23]),
     .sp4_v_b_07_16(net1112[0:47]), .sp4_h_l_07_16(net1068[0:47]),
     .slf_op_12_09(slf_op_12_09[7:0]),
     .bnl_op_12_09(slf_op_11_08[7:0]),
     .bot_op_12_09(slf_op_12_08[7:0]), .sp4_v_b_12_09(net727[0:47]),
     .sp12_v_b_12_09(net729[0:23]), .bnr_op_12_09({slf_op_13_08[3],
     slf_op_13_08[2], slf_op_13_08[1], slf_op_13_08[0],
     slf_op_13_08[3], slf_op_13_08[2], slf_op_13_08[1],
     slf_op_13_08[0]}), .slf_op_11_09(slf_op_11_09[7:0]),
     .bnl_op_11_09(slf_op_10_08[7:0]),
     .bot_op_11_09(slf_op_11_08[7:0]), .sp4_v_b_11_09(net733[0:47]),
     .sp12_v_b_11_09(net735[0:23]), .bnr_op_11_09(slf_op_12_08[7:0]),
     .slf_op_10_09(slf_op_10_09[7:0]),
     .bnl_op_10_09(slf_op_09_08[7:0]),
     .bot_op_10_09(slf_op_10_08[7:0]), .sp4_v_b_10_09(net739[0:47]),
     .sp12_v_b_10_09(net741[0:23]), .bnr_op_10_09(slf_op_11_08[7:0]),
     .slf_op_09_09(slf_op_09_09[7:0]),
     .bnl_op_09_09(slf_op_08_08[7:0]),
     .bot_op_09_09(slf_op_09_08[7:0]), .sp4_v_b_09_09(net745[0:47]),
     .sp12_v_b_09_09(net747[0:23]), .bnr_op_09_09(slf_op_10_08[7:0]),
     .slf_op_08_09(slf_op_08_09[7:0]),
     .bnl_op_08_09(slf_op_07_08[7:0]),
     .bot_op_08_09(slf_op_08_08[7:0]), .sp4_v_b_08_09(net751[0:47]),
     .sp12_v_b_08_09(net753[0:23]), .bnr_op_08_09(slf_op_09_08[7:0]),
     .lft_op_07_09(slf_op_06_09[7:0]),
     .slf_op_07_09(slf_op_07_09[7:0]), .sp12_h_l_07_09(net1081[0:23]),
     .sp4_v_b_07_09(net756[0:47]), .sp4_h_l_07_09(net1102[0:47]),
     .bot_op_07_09(slf_op_07_08[7:0]), .sp12_v_b_07_09(net758[0:23]),
     .bnr_op_07_09(slf_op_08_08[7:0]),
     .hold_t_r(fabric_out_08_17_ticegate),
     .hold_r_t(fabric_out_13_10_ricegate), .bm_sweb_i(bm_sweb_b2_o[1]),
     .bm_sdo_i(net974), .bm_sdi_i(bm_sdi_b2_o[1]),
     .bm_sclkrw_i(bm_sclkrw_b2_o[1]), .bm_sweb_o(net972),
     .bm_sdo_o(bm_sdo_b3_o), .bm_sdi_o(net974), .bm_sclkrw_o(net975),
     .update_i(net840), .tievdd(tievdd), .tiegnd(tiegnd),
     .tclk_i(tclkio_mr), .shift_i(net842), .sdi(sdio_mr), .r_i(net844),
     .purst(purst), .prog(prog), .mode_i(net845), .hiz_b_i(net846),
     .glb_in(gclk[7:0]), .ceb_i(net847), .bs_en_i(net848),
     .bm_wdummymux_en_i(net849), .bm_sreb_i(net851),
     .bm_sclk_i(net855), .bm_sa_i(net856[0:7]),
     .bm_rcapmux_en_i(net857), .bm_init_i(net858), .update_o(net1133),
     .tclk_o(tclkio_mt), .shift_o(net1137), .sdo(sdio_mt),
     .r_o(net1139), .mode_o(net1142), .hiz_b_o(net1143),
     .ceb_o(net1145), .bs_en_o(net1146), .bm_wdummymux_en_o(net1005),
     .bm_sreb_o(net1006), .bm_sclk_o(net1007), .bm_sa_o(net1008[0:7]),
     .bm_rcapmux_en_o(net1009), .bm_init_o(net1010));
ice1f_quad_tl I_quad_tl_ice1f ( .padin_l_t(padin_l[25:14]),
     .pado_l_t(pado_l[25:14]), .padeb_l_t(padeb_l[25:14]),
     .padeb_t_l(padeb_t[11:0]), .padin_t_l(padin_t[11:0]),
     .pado_t_l(pado_t[11:0]), .last_rsr(last_rsr),
     .carry_in_01_09(carry_io_01_0809),
     .carry_in_02_09(carry_io_02_0809),
     .carry_in_04_09(carry_io_04_0809),
     .carry_in_05_09(carry_io_05_0809),
     .carry_in_06_09(carry_io_06_0809), .sp12_v_b_06_09(net628[0:23]),
     .sp12_v_b_05_09(net552[0:23]), .bnr_op_05_09(slf_op_06_08[7:0]),
     .end_of_startup_top_l(end_of_startup_t[6:1]), .cf_t(cf_t[143:0]),
     .sp12_h_r_06_16(net1028[0:23]), .sp12_h_r_06_15(net1029[0:23]),
     .sp12_h_r_06_14(net1030[0:23]), .sp12_h_r_06_13(net1031[0:23]),
     .sp12_h_r_06_12(net1032[0:23]), .sp12_h_r_06_11(net1033[0:23]),
     .sp12_h_r_06_10(net1034[0:23]), .rgt_op_06_09(slf_op_07_09[7:0]),
     .fabric_out_00_09(fabric_out_00_09),
     .end_of_startup_lft_t(end_of_startup_l[16:9]),
     .sp12_v_b_01_09(net624[0:23]), .bot_op_05_09(slf_op_05_08[7:0]),
     .bot_op_04_09(slf_op_04_08[7:0]),
     .bot_op_03_09(slf_op_03_08[7:0]),
     .bot_op_02_09(slf_op_02_08[7:0]),
     .slf_op_02_09(slf_op_02_09[7:0]),
     .bnr_op_06_09(slf_op_07_08[7:0]),
     .bnr_op_04_09(slf_op_05_08[7:0]),
     .bnr_op_03_09(slf_op_04_08[7:0]),
     .bnr_op_02_09(slf_op_03_08[7:0]),
     .slf_op_00_09(slf_op_00_09[3:0]),
     .bnl_op_06_09(slf_op_05_08[7:0]),
     .bnl_op_05_09(slf_op_04_08[7:0]),
     .bnl_op_04_09(slf_op_03_08[7:0]),
     .bnl_op_03_09(slf_op_02_08[7:0]),
     .bnl_op_02_09(slf_op_01_08[7:0]),
     .bnr_op_01_09(slf_op_02_08[7:0]), .sp4_h_r_06_17(net1055[0:15]),
     .rgt_op_06_15(slf_op_07_15[7:0]),
     .rgt_op_06_14(slf_op_07_14[7:0]),
     .rgt_op_06_13(slf_op_07_13[7:0]),
     .rgt_op_06_12(slf_op_07_12[7:0]),
     .rgt_op_06_11(slf_op_07_11[7:0]),
     .rgt_op_06_10(slf_op_07_10[7:0]), .sp4_v_b_00_09(net598[0:15]),
     .bot_op_06_09(slf_op_06_08[7:0]),
     .slf_op_06_10(slf_op_06_10[7:0]),
     .slf_op_04_09(slf_op_04_09[7:0]),
     .rgt_op_06_16(slf_op_07_16[7:0]), .padin_00_09a(padin_0009a_ck),
     .sp4_h_r_06_16(net1068[0:47]), .bl(bl_top[329:0]),
     .vdd_cntl_l(vdd_cntl_l[287:144]),
     .bnr_op_00_09(slf_op_01_08[7:0]), .sp12_v_b_04_09(net627[0:23]),
     .sp12_v_b_03_09(net626[0:23]), .sp12_v_b_02_09(net625[0:23]),
     .sp4_r_v_b_06_15(net1075[0:47]), .sp4_r_v_b_06_14(net1076[0:47]),
     .sp4_r_v_b_06_13(net1077[0:47]), .sp4_r_v_b_06_12(net1078[0:47]),
     .sp4_r_v_b_06_11(net1079[0:47]), .sp4_r_v_b_06_10(net1080[0:47]),
     .sp12_h_r_06_09(net1081[0:23]), .bot_op_01_09(slf_op_01_08[7:0]),
     .sp4_v_b_06_09(net616[0:47]), .sp4_v_b_05_09(net615[0:47]),
     .sp4_v_b_04_09(net614[0:47]), .sp4_v_b_03_09(net613[0:47]),
     .sp4_v_b_02_09(net612[0:47]), .slf_op_01_09(slf_op_01_09[7:0]),
     .sp4_h_r_06_15(net1089[0:47]), .sp4_h_r_06_14(net1090[0:47]),
     .sp4_h_r_06_13(net1091[0:47]), .sp4_h_r_06_12(net1092[0:47]),
     .sp4_h_r_06_11(net1093[0:47]), .sp4_h_r_06_10(net1094[0:47]),
     .sp4_r_v_b_06_09(net756[0:47]), .slf_op_06_16(slf_op_06_16[7:0]),
     .slf_op_06_15(slf_op_06_15[7:0]),
     .slf_op_06_14(slf_op_06_14[7:0]),
     .slf_op_06_13(slf_op_06_13[7:0]),
     .slf_op_06_12(slf_op_06_12[7:0]),
     .slf_op_06_11(slf_op_06_11[7:0]), .sp4_h_r_06_09(net1102[0:47]),
     .reset_b_l(reset_b_l[287:144]), .pgate_l(pgate_l[287:144]),
     .fabric_out_06_17(fabric_out_06_17), .cf_l(cf_l[383:192]),
     .sp4_v_b_01_09(net611[0:47]), .tnr_op_06_16(slf_op_07_17[3:0]),
     .slf_op_06_09(slf_op_06_09[7:0]),
     .slf_op_05_09(slf_op_05_09[7:0]),
     .slf_op_03_09(slf_op_03_09[7:0]), .sp4_r_v_b_06_16(net1112[0:47]),
     .bnl_op_01_09({slf_op_00_08[3], slf_op_00_08[2], slf_op_00_08[1],
     slf_op_00_08[0], slf_op_00_08[3], slf_op_00_08[2],
     slf_op_00_08[1], slf_op_00_08[0]}),
     .slf_op_06_17(slf_op_06_17[3:0]), .padin_06_17b(padin_0617b_ck),
     .wl_l(wl_l[287:144]), .bm_init_o(bm_init_b1_o),
     .bm_sa_o(bm_sa_b1_o[7:0]), .bm_sclkrw_o(bm_sclkrw_b1_o),
     .bm_sclk_o(bm_sclk_b1_o), .bm_rcapmux_en_o(bm_rcapmux_en_b1_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_b1_o),
     .bm_sreb_o(bm_sreb_b1_o), .bm_sweb_o(bm_sweb_b1_o),
     .bm_sdi_o(bm_sdo_b1_i), .bm_sdo_i(bm_sdo_b1_i),
     .hold_t_l(fabric_out_08_17_ticegate),
     .hold_l_t(fabric_out_00_07_licegate), .bm_sweb_i(bm_sweb_b0_o[1]),
     .bm_sdi_i(bm_sdi_b0_o[1]), .bm_sclkrw_i(bm_sclkrw_b0_o[1]),
     .bm_sdo_o(bm_sdo_b1_o), .update_i(net1133), .tievdd(tievdd),
     .tiegnd(tiegnd), .tclk_i(tclkio_mt), .shift_i(net1137),
     .sdi(sdio_mt), .r_i(net1139), .purst(purst), .prog(prog),
     .mode_i(net1142), .hiz_b_i(net1143), .glb_in(gclk[7:0]),
     .ceb_i(net1145), .bs_en_i(net1146), .bm_wdummymux_en_i(net682),
     .bm_sreb_i(net684), .bm_sclk_i(net688), .bm_sa_i(net689[0:7]),
     .bm_rcapmux_en_i(net690), .bm_init_i(net691), .update_o(net649),
     .tclk_o(tclkio_ml), .shift_o(net653), .sdo(sdio_ml), .r_o(net655),
     .mode_o(net658), .hiz_b_o(net659), .ceb_o(net661),
     .bs_en_o(net662));
ice12p_clk_mux2to1 I_q4mux_ck5432 ( .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[145:144]), .bl(bl_top[333:330]),
     .min3({padin_1309a_ck, fabric_out_06_00}), .min2({padin_0009a_ck,
     fabric_out_06_17}), .min1({padin_0700a_ck, fabric_out_00_09}),
     .min0({padin_0717a_ck, fabric_out_13_09}), .wl_l(wl_l[145:144]),
     .reset_l(reset_b_l[145:144]), .pgate_l(pgate_l[145:144]),
     .gnet(gclk[5:2]), .pgate_r(pgate_r[145:144]),
     .wl_r(wl_r[145:144]), .reset_r(reset_b_r[145:144]),
     .vdd_cntl_r(vdd_cntl_r[145:144]));
ice12p_clk_mux2to1 I_q4mux_ck7610 ( .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[143:142]), .bl(bl_bot[333:330]),
     .min3({padin_0617b_ck, fabric_out_13_08}), .min2({padin_0600b_ck,
     fabric_out_00_08}), .min1({padin_0008b_ck, fabric_out_07_17}),
     .min0({padin_1308b_ck, fabric_out_07_00}), .wl_l(wl_l[143:142]),
     .reset_l(reset_b_l[143:142]), .pgate_l(pgate_l[143:142]),
     .gnet({gclk[7], gclk[6], gclk[1], gclk[0]}),
     .pgate_r(pgate_r[143:142]), .wl_r(wl_r[143:142]),
     .reset_r(reset_b_r[143:142]), .vdd_cntl_r(vdd_cntl_r[143:142]));
bram_bank_logic_bot I21 ( .bm_sdo_i(net852[0:1]),
     .bm_sclk_i(bm_bank30_sclk_o[1]), .bm_sclkrw_i(net1291),
     .bm_sweb_i(net1275), .bm_sdo_o(bm_bank30_sdo_i[3:2]),
     .bm_sweb_o(net831[0:1]), .bm_sclkrw_o(net835[0:1]),
     .bm_banksel_i(bm_bank30_banksel_o[3:2]));
bram_bank_logic_bot I10 ( .bm_sdo_i(net685[0:1]), .bm_sclk_i(net669),
     .bm_sclkrw_i(net1202), .bm_sweb_i(net1203),
     .bm_sdo_o(net1204[0:1]), .bm_sweb_o(net664[0:1]),
     .bm_sclkrw_o(net668[0:1]),
     .bm_banksel_i(bm_bank10_banksel_o[1:0]));
bram_hbuffer_2xbank I_bram_buf0 ( .bm_wdummymux_en_o(net1237),
     .bm_sweb_i(bm_sweb_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_init_i(bm_init_i), .bm_banksel_o(net1250[0:3]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_o(net1230),
     .bm_sreb_o(net1231), .bm_sclk_o(net1232), .bm_sa_o(net1233[0:7]),
     .bm_init_o(net1234), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclkrw_o(net1243), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sdo_o(bm_sdo_o[3:0]), .bm_sdi_o(net1245[0:3]),
     .bm_rcapmux_en_o(net1236), .bm_banksel_i(bm_banksel_i[3:0]),
     .bm_sdo_i(net1246[0:3]));
bram_hbuffer_dff_2xbank I_bram_buf1 ( .bm_sweb_i(net1230),
     .bm_sreb_i(net1231), .bm_sclk_i(net1232), .bm_sa_i(net1233[0:7]),
     .bm_init_i(net1234), .bm_banksel_o(bm_bank30_banksel_o[3:0]),
     .bm_rcapmux_en_i(net1236), .bm_wdummymux_en_i(net1237),
     .bm_sweb_o(net1275), .bm_sreb_o(net1276),
     .bm_sclk_o(bm_bank30_sclk_o[1:0]), .bm_sa_o(net1279[0:7]),
     .bm_init_o(net1280), .bm_sclkrw_i(net1243), .bm_sclkrw_o(net1291),
     .bm_sdi_i(net1245[0:3]), .bm_sdo_o(net1246[0:3]),
     .bm_sdi_o(bm_bank30_sdi_o[3:0]), .bm_rcapmux_en_o(net1282),
     .bm_wdummymux_en_o(net1283), .bm_banksel_i(net1250[0:3]),
     .bm_sdo_i(bm_bank30_sdo_i[3:0]));
bram_hbuffer_1xbank I_bram_buf3 ( .bm_wdummymux_en_o(net663),
     .bm_sweb_i(net1253), .bm_sreb_i(net1254), .bm_sdi_i(net1255[0:1]),
     .bm_sclk_i(net1256), .bm_sa_i(net1257[0:7]), .bm_init_i(net1258),
     .bm_banksel_o(bm_bank10_banksel_o[1:0]),
     .bm_rcapmux_en_i(net1260), .bm_wdummymux_en_i(net1261),
     .bm_sweb_o(net1203), .bm_sreb_o(net665), .bm_sdi_o(net667[0:1]),
     .bm_sclk_o(net669), .bm_sa_o(net670[0:7]), .bm_init_o(net672),
     .bm_rcapmux_en_o(net671), .bm_sclkrw_i(net1269),
     .bm_sclkrw_o(net1202), .bm_sdo_i(net1204[0:1]),
     .bm_banksel_i(net1272[0:1]), .bm_sdo_o(net1273[0:1]));
bram_hbuffer_1xbank I_bram_buf2 ( .bm_wdummymux_en_o(net1261),
     .bm_sweb_i(net1275), .bm_sreb_i(net1276),
     .bm_sdi_i(bm_bank30_sdi_o[1:0]), .bm_sclk_i(bm_bank30_sclk_o[0]),
     .bm_sa_i(net1279[0:7]), .bm_init_i(net1280),
     .bm_banksel_o(net1272[0:1]), .bm_rcapmux_en_i(net1282),
     .bm_wdummymux_en_i(net1283), .bm_sweb_o(net1253),
     .bm_sreb_o(net1254), .bm_sdi_o(net1255[0:1]), .bm_sclk_o(net1256),
     .bm_sa_o(net1257[0:7]), .bm_init_o(net1258),
     .bm_rcapmux_en_o(net1260), .bm_sclkrw_i(net1291),
     .bm_sclkrw_o(net1269), .bm_sdo_i(net1273[0:1]),
     .bm_banksel_i(bm_bank30_banksel_o[1:0]),
     .bm_sdo_o(bm_bank30_sdo_i[1:0]));

endmodule
// Library - leafcell, Cell - tielo4x, View - schematic
// LAST TIME SAVED: Sep 10 09:05:31 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module tielo4x ( tielo );
output  tielo;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M0 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));
nch_hvt  M1 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - leafcell, Cell - tiehi4x, View - schematic
// LAST TIME SAVED: Sep 10 09:03:54 2007
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module tiehi4x ( tiehi );
output  tiehi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - chip, Cell - chip_ice1f, View - schematic
// LAST TIME SAVED: Jul 20 12:19:11 2009
// NETLIST TIME: Aug 24 09:59:03 2009
`timescale 1ns / 1ns 

module chip_ice1f ( tdo, cdone, uio_bbank, uio_lbank, uio_rbank,
     uio_tbank, vpp, creset_b, tck, tdi, tms, trstb );

output  tdo;

inout  cdone, vpp;

input  creset_b, tck, tdi, tms, trstb;

inout [25:0]  uio_lbank;
inout [23:0]  uio_bbank;
inout [20:0]  uio_rbank;
inout [23:0]  uio_tbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net135;

wire  [3:0]  bm_sdo_o;

wire  [23:12]  spi_ss_in_bbank;

wire  [287:0]  pgate_r;

wire  [31:0]  spi_ss_in_r;

wire  [663:0]  bl_top;

wire  [287:0]  cf_tbank;

wire  [287:0]  reset_l;

wire  [25:0]  out_lbank;

wire  [287:0]  wl_l;

wire  [287:0]  reset_r;

wire  [25:0]  in_lbank;

wire  [20:0]  oen_rbank;

wire  [23:0]  oen_tbank;

wire  [383:0]  cf_lbank;

wire  [287:0]  wl_r;

wire  [3:0]  bm_sdi_o;

wire  [23:0]  out_tbank;

wire  [23:0]  oen_bbank;

wire  [287:0]  vdd_cntl_l;

wire  [23:0]  in_tbank;

wire  [287:0]  vdd_cntl_r;

wire  [287:0]  cf_bbank;

wire  [20:0]  out_rbank;

wire  [20:0]  in_rbank;

wire  [25:0]  oen_lbank;

wire  [663:0]  bl_bot;

wire  [3:0]  bm_banksel_i;

wire  [23:0]  in_bbank;

wire  [23:0]  out_bbank;

wire  [3:0]  last_rsr;

wire  [383:0]  cf_rbank;

wire  [7:0]  bm_sa_i;

wire  [287:0]  pgate_l;

wire  [0:6]  net131;



ring_route_ice1f_july16 I_ring_route1f ( .out_rbank(out_rbank[20:0]),
     .out_bbank({out_bbank[23:13], out_bbank[11], out_bbank[10],
     out_bbank[12], out_bbank[9:0]}), .oen_rbank(oen_rbank[20:0]),
     .oen_bbank({oen_bbank[23:13], oen_bbank[11], oen_bbank[10],
     oen_bbank[12], oen_bbank[9:0]}), .cf_rbank({cf_rbank[346],
     cf_rbank[336], cf_rbank[322], cf_rbank[312], cf_rbank[298],
     cf_rbank[288], cf_rbank[274], cf_rbank[264], cf_rbank[250],
     cf_rbank[240], cf_rbank[202], cf_rbank[192], cf_rbank[178],
     cf_rbank[168], cf_rbank[154], cf_rbank[144], cf_rbank[130],
     cf_rbank[120], cf_rbank[82], cf_rbank[72], cf_rbank[58]}),
     .cf_bbank({cf_bbank[274], cf_bbank[264], cf_bbank[250],
     cf_bbank[240], cf_bbank[226], cf_bbank[216], cf_bbank[202],
     cf_bbank[192], cf_bbank[178], cf_bbank[168], cf_bbank[154],
     cf_bbank[130], cf_bbank[120], cf_bbank[144], cf_bbank[106],
     cf_bbank[96], cf_bbank[82], cf_bbank[72], cf_bbank[58],
     cf_bbank[48], cf_bbank[34], cf_bbank[24], cf_bbank[10],
     cf_bbank[0]}), .in_rbank(in_rbank[20:0]),
     .in_bbank({in_bbank[23:13], in_bbank[11], in_bbank[10],
     in_bbank[12], in_bbank[9:0]}), .uio_rbank(uio_rbank[20:0]),
     .uio_bbank(uio_bbank[23:0]), .uio_lbank(uio_lbank[25:0]),
     .in_lbank(in_lbank[25:0]), .cf_lbank({cf_lbank[383], cf_lbank[23],
     cf_lbank[322], cf_lbank[312], cf_lbank[298], cf_lbank[288],
     cf_lbank[274], cf_lbank[264], cf_lbank[250], cf_lbank[240],
     cf_lbank[226], cf_lbank[216], cf_lbank[202], cf_lbank[192],
     cf_lbank[178], cf_lbank[168], cf_lbank[130], cf_lbank[120],
     cf_lbank[106], cf_lbank[96], cf_lbank[82], cf_lbank[72],
     cf_lbank[58], cf_lbank[48], cf_lbank[34], cf_lbank[24],
     cf_lbank[10], cf_lbank[0]}), .oen_lbank(oen_lbank[25:0]),
     .out_lbank(out_lbank[25:0]), .uio_tbank(uio_tbank[23:0]),
     .in_tbank(in_tbank[23:0]), .oen_tbank(oen_tbank[23:0]),
     .out_tbank(out_tbank[23:0]), .cf_tbank({cf_tbank[274],
     cf_tbank[264], cf_tbank[250], cf_tbank[240], cf_tbank[226],
     cf_tbank[216], cf_tbank[202], cf_tbank[192], cf_tbank[178],
     cf_tbank[168], cf_tbank[154], cf_tbank[144], cf_tbank[130],
     cf_tbank[120], cf_tbank[106], cf_tbank[96], cf_tbank[82],
     cf_tbank[72], cf_tbank[58], cf_tbank[48], cf_tbank[34],
     cf_tbank[24], cf_tbank[10], cf_tbank[0]}),
     .spi_ss_in_bbank(spi_ss_in_bbank[23:18]), .en_8bconfig_b(net130),
     .psdo(net131[0:6]), .fabric_out_12_00(wb_boot),
     .fabric_out_13_01(wb_boot_sel0), .fabric_out_13_02(wb_boot_sel1),
     .trstb(trstb), .tms(tms), .tdi(tdi), .tck(tck),
     .spi_ss_in_r({tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd}), .fromsdo(fromsdo), .creset_b(creset_b),
     .bm_sdo_o(bm_sdo_o[3:0]), .vdd_cntl_r(vdd_cntl_r[287:0]),
     .vdd_cntl_l(vdd_cntl_l[287:0]), .update0(update0), .tdo(tdo),
     .j_tck(j_tck), .spi_ss_out_b(spi_ss_out_b),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .spi_clk_out(spi_clk_out), .shift0(shift0),
     .reset_r(reset_r[287:0]), .reset_l(reset_l[287:0]),
     .pgate_r(pgate_r[287:0]), .pgate_l(pgate_l[287:0]), .mode0(mode0),
     .md_spi_b(md_spi_b), .last_rsr(last_rsr[3:0]),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .j_tdi(j_tdi), .hiz_b0(hiz_b0), .gsr(gsr), .gint_hz(gint_hz),
     .end_of_startup(end_of_startup), .bs_en0(bs_en0),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sdi_i(bm_sdi_o[3:0]),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .bm_banksel_i(bm_banksel_i[3:0]),
     .cdone(cdone), .bl_top(bl_top[663:0]), .bl_bot(bl_bot[663:0]),
     .cf_r_ext({cf_rbank[383], cf_rbank[23]}), .tiegnd(tiegnd),
     .tievdd(tievdd), .vpp(vpp), .ceb0(ceb), .wl_l(wl_l[287:0]),
     .wl_r(wl_r[287:0]));
ice1f_quad_x4 I_ICE1f_quad_x4 ( .padeb_b(oen_bbank[23:0]),
     .pado_b(out_bbank[23:0]), .padin_b(in_bbank[23:0]),
     .padeb_r(oen_rbank[20:0]), .pado_r(out_rbank[20:0]),
     .padin_r(in_rbank[20:0]), .padeb_l(oen_lbank[25:0]),
     .pado_l(out_lbank[25:0]), .padin_l(in_lbank[25:0]),
     .pado_t(out_tbank[23:0]), .padeb_t(oen_tbank[23:0]),
     .padin_t(in_tbank[23:0]), .last_rsr(last_rsr[1]),
     .end_of_startup_b({end_of_startup, end_of_startup, end_of_startup,
     tievdd, tievdd, tievdd}), .vdd_cntl_r(vdd_cntl_r[287:0]),
     .vdd_cntl_l(vdd_cntl_l[287:0]), .update(update0), .tievdd(tievdd),
     .tiegnd(tiegnd), .tclk(j_tck), .spiout_r({tiegnd, tiegnd, tiegnd,
     last_rsr[3], tiegnd, last_rsr[2], tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .spiout_l({tiegnd, last_rsr[0], tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd}), .spioeb_l({tievdd, tiegnd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd}), .shift(shift0), .sdi_pad(j_tdi),
     .reset_b_r(reset_r[287:0]), .reset_b_l(reset_l[287:0]), .r(gsr),
     .purst(gsr), .prog(gint_hz), .pgate_r(pgate_r[287:0]),
     .pgate_l(pgate_l[287:0]), .mode(mode0), .hiz_b(hiz_b0),
     .end_of_startup_t({tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}),
     .end_of_startup_r({tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, jtag_rowtest_mode_rowu3_b,
     jtag_rowtest_mode_rowu2_b, tievdd, tievdd, tievdd, tievdd,
     tievdd}), .end_of_startup_l({tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu0_b, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd}), .ceb(ceb), .bs_en(bs_en0),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sdi_i(bm_sdi_o[3:0]),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .bm_banksel_i(bm_banksel_i[3:0]),
     .spi_ss_in_r(spi_ss_in_r[31:0]), .spi_ss_in_l(net135[0:15]),
     .sdo_pad(fromsdo), .fabric_out_13_01_wb_sel0(wb_boot_sel0),
     .bm_sdo_o(bm_sdo_o[3:0]), .wl_l(wl_l[287:0]),
     .cf_l(cf_lbank[383:0]), .cf_b(cf_bbank[287:0]),
     .bl_top(bl_top[663:0]), .bl_bot(bl_bot[663:0]),
     .fabric_out_12_00_wb(wb_boot), .wl_r(wl_r[287:0]),
     .cf_t(cf_tbank[287:0]), .cf_r(cf_rbank[383:0]),
     .fabric_out_13_02_wb_sel1(wb_boot_sel1), .spiout_b({spi_ss_out_b,
     spi_clk_out, tiegnd, spi_sdo, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd}), .spioeb_b({md_spi_b, md_spi_b,
     tievdd, spi_sdo_oe_b, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd}), .spi_ss_in_b(spi_ss_in_bbank[23:12]));
tielo4x I_tielo ( .tielo(tiegnd));
tiehi4x I_tiehi ( .tiehi(tievdd));

endmodule
// Library - misc, Cell - ml_osc_top, View - schematic
// LAST TIME SAVED: Oct 14 15:44:25 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_osc_top ( cnt_podt_out, smc_clk, crst_b, por_b, smc_osc_fsel,
     smc_oscoff_b, smc_podt_off, smc_podt_rst );
output  cnt_podt_out, smc_clk;

input  crst_b, por_b, smc_oscoff_b, smc_podt_off, smc_podt_rst;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:0]  q_b;

wire  [10:0]  q;



tiehi I179 ( .tiehi(net076));
nor2_hvt I256 ( .A(rst_osc_b), .B(smc_oscoff_b), .Y(net066));
nor2_hvt I266 ( .A(clk_out), .B(smc_podt_off), .Y(net078));
nor2_hvt I257 ( .A(disable_osc), .B(net066), .Y(smc_oscen));
nor2_hvt I264 ( .A(smc_podt_rst), .B(net090), .Y(net054));
nor2_hvt I252 ( .A(cnt_rst), .B(smc_oscoff_b), .Y(net0124));
nand2_hvt I227 ( .A(smc_off_b), .B(rst_osc_b), .Y(disable_osc));
nand2_hvt I270 ( .A(crst_b), .Y(net064), .B(por_b));
ml_dff I230 ( .R(cnt_rst), .D(net076), .CLK(q_b[10]), .QN(net067),
     .Q(net063));
ml_dff I243 ( .R(rst_off_latch), .D(net0174), .CLK(clk_out_b),
     .QN(smc_off_b), .Q(net0152));
ml_dff I228_10_ ( .R(cnt_rst), .D(q_b[10]), .CLK(q[9]), .QN(q_b[10]),
     .Q(q[10]));
ml_dff I228_9_ ( .R(cnt_rst), .D(q_b[9]), .CLK(q[8]), .QN(q_b[9]),
     .Q(q[9]));
ml_dff I228_8_ ( .R(cnt_rst), .D(q_b[8]), .CLK(q[7]), .QN(q_b[8]),
     .Q(q[8]));
ml_dff I228_7_ ( .R(cnt_rst), .D(q_b[7]), .CLK(q[6]), .QN(q_b[7]),
     .Q(q[7]));
ml_dff I228_6_ ( .R(cnt_rst), .D(q_b[6]), .CLK(q[5]), .QN(q_b[6]),
     .Q(q[6]));
ml_dff I228_5_ ( .R(cnt_rst), .D(q_b[5]), .CLK(q[4]), .QN(q_b[5]),
     .Q(q[5]));
ml_dff I228_4_ ( .R(cnt_rst), .D(q_b[4]), .CLK(q[3]), .QN(q_b[4]),
     .Q(q[4]));
ml_dff I228_3_ ( .R(cnt_rst), .D(q_b[3]), .CLK(q[2]), .QN(q_b[3]),
     .Q(q[3]));
ml_dff I228_2_ ( .R(cnt_rst), .D(q_b[2]), .CLK(q[1]), .QN(q_b[2]),
     .Q(q[2]));
ml_dff I228_1_ ( .R(cnt_rst), .D(q_b[1]), .CLK(q[0]), .QN(q_b[1]),
     .Q(q[1]));
ml_dff I228_0_ ( .R(cnt_rst), .D(q_b[0]), .CLK(clk_in), .QN(q_b[0]),
     .Q(q[0]));
inv_hvt I233 ( .A(clk_out), .Y(clk_out_b));
inv_hvt I271 ( .A(net064), .Y(rst_osc_b));
inv_hvt I267 ( .A(net078), .Y(clk_in));
inv_hvt I262 ( .A(net067), .Y(cnt_podt_out));
inv_hvt I244 ( .A(smc_oscoff_b), .Y(net0174));
inv_hvt I265 ( .A(net054), .Y(cnt_rst));
inv_hvt I229 ( .A(rst_osc_b), .Y(net090));
inv_hvt I253 ( .A(net0124), .Y(rst_off_latch));
inv_hvt I232 ( .A(clk_out_b), .Y(smc_clk));
ml_osc Iml_osc ( .smc_osc_fsel(smc_osc_fsel[1:0]), .clk_out(clk_out),
     .smc_oscen(smc_oscen));

endmodule
// Library - leafcell, Cell - bram_bufferx16, View - schematic
// LAST TIME SAVED: Jun 25 13:49:31 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module bram_bufferx16 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I0 ( .A(net07), .Y(net09));
inv_hvt I2 ( .A(in), .Y(net07));
inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(net09), .Y(net6));

endmodule
// Library - xpmem, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jun  5 11:34:46 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - xpmem, Cell - ml_cram_logic, View - schematic
// LAST TIME SAVED: Sep 28 20:58:40 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_cram_logic ( cram_pgateoff, cram_prec, cram_pullup_b,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, smc_clk_out, por,
     smc_clk, smc_read, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rwl_en, smc_seq_rst, smc_wcram_rst, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en );
output  cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, smc_clk_out;

input  por, smc_clk, smc_read, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_write, smc_wset_prec, smc_wset_precgnd, smc_wwlwrt_dis,
     smc_wwlwrt_en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I213 ( .A(net208), .Y(net177), .B(net248));
inv_hvt I370 ( .A(net273), .Y(rst_rpull_rwl));
inv_hvt I373 ( .A(cram_rst), .Y(net257));
inv_hvt I346 ( .A(net315), .Y(net220));
inv_hvt I263 ( .A(net269), .Y(net218));
inv_hvt I266 ( .A(cram_write_int), .Y(net216));
inv_hvt I286 ( .A(net359), .Y(net299));
inv_hvt I422 ( .A(smc_rwl_en), .Y(net212));
inv_hvt I323 ( .A(net282), .Y(net210));
inv_hvt I378 ( .A(net276), .Y(net248));
inv_hvt I333 ( .A(net279), .Y(net208));
inv_hvt I324 ( .A(net210), .Y(cram_pgateoff));
inv_hvt I403 ( .A(net285), .Y(net204));
inv_hvt I292 ( .A(net200), .Y(cram_prec));
inv_hvt I267 ( .A(net303), .Y(net200));
inv_hvt I224 ( .A(net291), .Y(reset_logic));
inv_hvt I401 ( .A(net294), .Y(net196));
inv_hvt I381 ( .A(net309), .Y(net194));
inv_hvt I268 ( .A(net257), .Y(net253));
inv_hvt I293 ( .A(net236), .Y(cram_vddoff));
inv_hvt I269 ( .A(net255), .Y(net251));
inv_hvt I330 ( .A(net265), .Y(net190));
inv_hvt I374 ( .A(net253), .Y(net255));
inv_hvt I294 ( .A(cram_rst_int_b), .Y(cram_rst));
inv_hvt I375 ( .A(net252), .Y(cram_rst_dly));
inv_hvt I421 ( .A(net394), .Y(net186));
inv_hvt I249 ( .A(net262), .Y(net184));
inv_hvt I250 ( .A(net184), .Y(cram_pullup_b));
inv_hvt I359 ( .A(net179), .Y(net180));
inv_hvt I376 ( .A(net251), .Y(net252));
inv_hvt I336 ( .A(smc_clk), .Y(sm_clk_b));
inv_hvt I367 ( .A(net306), .Y(dis_pgatewrt));
inv_hvt I281 ( .A(net399), .Y(net226));
inv_hvt I399 ( .A(net300), .Y(net240));
inv_hvt I290 ( .A(net218), .Y(cram_wl_en));
inv_hvt I425 ( .A(net299), .Y(net262));
inv_hvt I337 ( .A(sm_clk_b), .Y(smc_clk_out));
inv_hvt I256 ( .A(net379), .Y(cram_write_int));
inv_hvt I291 ( .A(net216), .Y(cram_write));
inv_hvt I415 ( .A(net312), .Y(net260));
inv_hvt I312 ( .A(net177), .Y(net228));
inv_hvt I270 ( .A(net228), .Y(net236));
inv_hvt I271 ( .A(net226), .Y(cram_rst_int_b));
mux2_hvt I161 ( .in1(cram_write_int), .in0(net186), .out(net269),
     .sel(net208));
mux2_hvt I295 ( .in1(net194), .in0(net220), .out(net265),
     .sel(net208));
nor2_hvt I402 ( .A(net283), .B(smc_wset_precgnd), .Y(net285));
nor2_hvt I329 ( .A(net190), .B(smc_seq_rst), .Y(net303));
nor2_hvt I398 ( .A(smc_rpull_b), .B(net299), .Y(net300));
nor2_hvt I393 ( .A(cram_rst_dly), .B(reset_logic), .Y(net179));
nor2_hvt I364 ( .A(net389), .B(smc_seq_rst), .Y(net282));
nor2_hvt I400 ( .A(net292), .B(smc_wset_prec), .Y(net294));
nor2_hvt I366 ( .A(reset_logic), .B(net370), .Y(net306));
nor2_hvt I223 ( .A(net318), .B(por), .Y(net291));
nor2_hvt I390 ( .A(smc_write), .B(smc_seq_rst), .Y(net279));
nor2_hvt I392 ( .A(net283), .B(cram_rst), .Y(net276));
nor2_hvt I389 ( .A(net375), .B(reset_logic), .Y(net273));
nor2_hvt I385 ( .A(smc_rprec), .B(net287), .Y(net315));
nor2_hvt I414 ( .A(net310), .B(smc_wwlwrt_en), .Y(net312));
nor2_hvt I391 ( .A(net292), .B(cram_rst), .Y(net309));
nor3_hvt I220 ( .B(net322), .Y(net326), .A(net322), .C(net322));
nor3_hvt I217 ( .B(net401), .Y(net330), .A(net401), .C(net401));
nor3_hvt I386 ( .B(smc_seq_rst), .Y(net318), .A(smc_write),
     .C(smc_read));
nor3_hvt I218 ( .B(net330), .Y(net322), .A(net330), .C(net330));
nor3_hvt I387 ( .B(smc_rwl_en), .Y(net287), .A(net315),
     .C(reset_logic));
nand3_hvt I230 ( .Y(net348), .B(net344), .C(net344), .A(net344));
nand3_hvt I231 ( .Y(net352), .B(net348), .C(net348), .A(net348));
nand3_hvt I426 ( .Y(net344), .B(net401), .C(net401), .A(net401));
ml_dff_schematic I411 ( .R(reset_logic), .D(smc_wwlwrt_dis),
     .CLK(smc_clk), .QN(net369), .Q(net370));
ml_dff_schematic I408 ( .R(rst_rpull_rwl), .D(net401), .CLK(net212),
     .QN(net394), .Q(net395));
ml_dff_schematic I405 ( .R(dis_pgatewrt), .D(net401),
     .CLK(cram_rst_int_b), .QN(net389), .Q(net390));
ml_dff_schematic I412 ( .R(net180), .D(net196), .CLK(smc_clk_out),
     .QN(net337), .Q(net292));
ml_dff_schematic I410 ( .R(dis_pgatewrt), .D(net260),
     .CLK(smc_clk_out), .QN(net379), .Q(net310));
ml_dff_schematic I108 ( .R(reset_logic), .D(smc_rrst_pullwlen),
     .CLK(smc_clk_out), .QN(net343), .Q(net375));
ml_dff_schematic I413 ( .R(net180), .D(net204), .CLK(smc_clk_out),
     .QN(net333), .Q(net283));
ml_dff_schematic I407 ( .R(rst_rpull_rwl), .D(net240),
     .CLK(smc_clk_out), .QN(net359), .Q(net360));
ml_dff_schematic I406 ( .R(reset_logic), .D(smc_wcram_rst),
     .CLK(smc_clk_out), .QN(net399), .Q(net400));
tiehi I427 ( .tiehi(net401));

endmodule
// Library - chip, Cell - CHIP_smc_ice12k, View - schematic
// LAST TIME SAVED: Aug 14 11:21:37 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module CHIP_smc_ice12k ( bm_banksel_i, bm_init_i, bm_rcapmux_en_i,
     bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bs_en0, cdone_out, ceb0, cm_banksel,
     cm_banksel_blbrd_2_, cm_banksel_bldld, cm_sdi_u0, cm_sdi_u1,
     cm_sdi_u2d, cm_sdi_u3, core_por_b0, core_por_bb, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, data_muxsel, data_muxsel1, en_8bconfig_b,
     end_of_startup, gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     md_spi_b, mode0, nvcm_spi_sdi, nvcm_spi_ss_b, psdo, row_test0,
     rst_b, sdo_enable, shift0, smc_clk_out, smc_load_nvcm_bstream,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk, smc_write0, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out_b, totdopad, update0, bm_sdo_o,
     bp0, cdone_in, cm_sdo_u0d1, cm_sdo_u1d3, cm_sdo_u2d1, cm_sdo_u3d1,
     creset_b_int, fabric_out_40_00, fabric_out_41_01,
     fabric_out_41_02, fromsdo, idcode_msb20bits, last_rsr3,
     monitor_celld4, monitor_celld, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, spi_ss_in_bbank,
     spi_ss_in_r, tck_pad, tdi_pad, tms_pad, trst_pad, vddio_rightbank
     );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, core_por_b0, core_por_bb, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, data_muxsel, data_muxsel1, en_8bconfig_b,
     end_of_startup, gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     md_spi_b, mode0, nvcm_spi_sdi, nvcm_spi_ss_b, row_test0, rst_b,
     sdo_enable, shift0, smc_clk_out, smc_load_nvcm_bstream,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk, smc_write0, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out_b, totdopad, update0;

input  bp0, cdone_in, creset_b_int, fabric_out_40_00, fabric_out_41_01,
     fabric_out_41_02, fromsdo, last_rsr3, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, tck_pad, tdi_pad,
     tms_pad, trst_pad, vddio_rightbank;

output [1:0]  cm_sdi_u1;
output [1:0]  cm_banksel_bldld;
output [3:0]  bm_sdi_i;
output [3:0]  bm_banksel_i;
output [1:0]  cm_sdi_u2d;
output [7:0]  bm_sa_i;
output [1:0]  cm_sdi_u3;
output [3:0]  cm_banksel;
output [7:1]  psdo;
output [1:0]  cm_sdi_u0;

input [1:0]  cm_sdo_u0d1;
input [4:0]  spi_ss_in_bbank;
input [19:0]  idcode_msb20bits;
input [1:0]  cm_sdo_u1d3;
input [7:1]  spi_ss_in_r;
input [1:0]  monitor_celld4;
input [3:2]  monitor_celld;
input [1:0]  cm_sdo_u2d1;
input [3:0]  bm_sdo_o;
input [1:0]  cm_sdo_u3d1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:1]  spi_ss_in_rd;

wire  [1:0]  u1_in;

wire  [1:0]  u0_in;

wire  [4:0]  spi_ss_in_bbankd;

wire  [1:0]  cm_sdi_u2;

wire  [1:0]  smc_osco_fsel;



creset_filter I14 ( .in(creset_b_int), .out(crst_filterout));
fabric_buf8k I1 ( .f_in(net281), .f_out(gsr));
fabric_buf8k I2 ( .f_in(net282), .f_out(gint_hz));
fabric_buf8k I3 ( .f_in(net283), .f_out(end_of_startup));
smc_and_jtag I_smc_and_jtag ( .warmboot_sel({fabric_out_41_02,
     fabric_out_41_01}), .trst_pad(trst_pad), .tms_pad(tms_pad),
     .tdi_pad(tdi_pad), .tck_pad(tck_pad),
     .spi_ss_in_b(spi_ss_in_bbankd[4]), .cnt_podt_out(cnt_podt_out),
     .spi_sdi(spi_ss_in_bbankd[2]), .spi_clk_in(spi_ss_in_bbankd[3]),
     .psdi(spi_ss_in_rd[7:1]), .por_b(smc_por_b0), .osc_clk(osc_clk),
     .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_spi_sdo(nvcm_spi_sdo), .nvcm_relextspi(nvcm_relextspi),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot),
     .creset_b(crst_filterout), .coldboot_sel(spi_ss_in_bbankd[1:0]),
     .cm_sdo_u2(cm_sdo_u2d1[1:0]), .cm_sdo_u1(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0(cm_sdo_u0d1[1:0]), .cm_sdi_u3(cm_sdi_u3[1:0]),
     .cm_monitor_cell({monitor_celld[3:2], monitor_celld4[1:0]}),
     .cm_last_rsr(last_rsr3), .cdone_in(cdone_in),
     .bschain_sdo(fromsdo), .bp0(bp0), .boot(fabric_out_40_00),
     .bm_bank_sdo(bm_sdo_o[3:0]), .tdo_pad(totdopad),
     .tdo_oe_pad(sdo_enable), .spi_ss_out_b(spi_ss_out_b),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .spi_clk_out(spi_clk_outd), .smc_wwlwrt_en(net246),
     .smc_wwlwrt_dis(net247), .smc_wset_precgnd(net248),
     .smc_wset_prec(net249), .smc_write(smc_write),
     .smc_wdis_dclk(smc_wdis_dclkd), .smc_wcram_rst(net252),
     .smc_seq_rst(net253), .smc_rwl_en(net254),
     .smc_rsr_rst(smc_rsr_rstd), .smc_rrst_pullwlen(net256),
     .smc_rpull_b(net257), .smc_rprec(net258),
     .smc_row_inc(smc_row_incd), .smc_read(net260),
     .smc_podt_rst(smc_podt_rst), .smc_podt_off(smc_podt_off),
     .smc_oscoff_b(smc_oscoff_b), .smc_osc_fsel(smc_osco_fsel[1:0]),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .psdo(psdo[7:1]), .nvcm_spi_ss_b(nvcm_spi_ss_b),
     .nvcm_spi_sdi(nvcm_spi_sdi), .md_spi_b(md_spi_b),
     .j_upd_dr(update0), .j_tdi(j_tdi), .j_tck(net0272),
     .j_shift0(shift0), .j_sft_dr(shiftfromsmc), .j_rst_b(j_rst_b),
     .j_row_test(row_test0), .j_mode(mode0), .j_hiz_b(hiz_b0),
     .j_ceb0(ceb0), .gsr(net281), .gint_hz(net282),
     .end_of_startup(net283), .en_8bconfig_b(en_8bconfig_b),
     .data_muxsel1(data_muxsel1d), .data_muxsel(data_muxseld),
     .cm_sdi_u2(cm_sdi_u2[1:0]), .cm_sdi_u1(u1_in[1:0]),
     .cm_sdi_u0(u0_in[1:0]), .cm_clk(net290),
     .cm_banksel(cm_banksel[3:0]), .cdone_out(cdone_out),
     .bs_en(bs_en0), .bm_wdummymux_en(bm_wdummymux_en_i),
     .bm_sweb(bm_sweb_i), .bm_sreb(bm_sreb_i), .bm_sclkrw(bm_sclkrw_i),
     .bm_sa(bm_sa_i[7:0]), .bm_rcapmux_en(bm_rcapmux_en_i),
     .bm_init(bm_init_i), .bm_clk(bm_sclk_i),
     .bm_banksel(bm_banksel_i[3:0]), .bm_bank_sdi(bm_sdi_i[3:0]),
     .idcode_msb20bits(idcode_msb20bits[19:0]),
     .cm_sdo_u3(cm_sdo_u3d1[1:0]));
SMC_CORE_POR_right I11 ( .creset_b(crst_filterout),
     .vddio_rightbank(vddio_rightbank), .smc_por_b(smc_por_b0),
     .core_por_b(core_por_b0),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2));
sg_bufx10 I15 ( .in(data_muxseld), .out(data_muxsel));
sg_bufx10 I16 ( .in(data_muxsel1d), .out(data_muxsel1));
sg_bufx10 I21 ( .in(net0272), .out(j_tck));
sg_bufx10 I18 ( .in(smc_rsr_rstd), .out(smc_rsr_rst));
sg_bufx10 I17 ( .in(smc_write), .out(smc_write0));
sg_bufx10 I19 ( .in(smc_row_incd), .out(smc_row_inc));
sg_bufx10 I5 ( .in(smc_wdis_dclkd), .out(smc_wdis_dclk));
sg_bufx10 I4_1_ ( .in(u1_in[1]), .out(cm_sdi_u1[1]));
sg_bufx10 I4_0_ ( .in(u1_in[0]), .out(cm_sdi_u1[0]));
sg_bufx10 I9_1_ ( .in(cm_sdi_u2[1]), .out(cm_sdi_u2d[1]));
sg_bufx10 I9_0_ ( .in(cm_sdi_u2[0]), .out(cm_sdi_u2d[0]));
sg_bufx10 I6_1_ ( .in(u0_in[1]), .out(cm_sdi_u0[1]));
sg_bufx10 I6_0_ ( .in(u0_in[0]), .out(cm_sdi_u0[0]));
sg_bufx10 I10 ( .in(cm_banksel[2]), .out(cm_banksel_blbrd_2_));
sg_bufx10 I13_1_ ( .in(cm_banksel[1]), .out(cm_banksel_bldld[1]));
sg_bufx10 I13_0_ ( .in(cm_banksel[0]), .out(cm_banksel_bldld[0]));
sg_bufx10 I0 ( .in(spi_clk_outd), .out(spi_clk_out));
inv_hvt I12 ( .A(core_por_b0), .Y(core_por_bb));
ml_osc_top Iml_osc ( .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]), .por_b(core_por_b0),
     .crst_b(crst_filterout), .smc_clk(osc_clk),
     .cnt_podt_out(cnt_podt_out));
bram_bufferx16 I20_4_ ( .in(spi_ss_in_bbank[4]),
     .out(spi_ss_in_bbankd[4]));
bram_bufferx16 I20_3_ ( .in(spi_ss_in_bbank[3]),
     .out(spi_ss_in_bbankd[3]));
bram_bufferx16 I20_2_ ( .in(spi_ss_in_bbank[2]),
     .out(spi_ss_in_bbankd[2]));
bram_bufferx16 I20_1_ ( .in(spi_ss_in_bbank[1]),
     .out(spi_ss_in_bbankd[1]));
bram_bufferx16 I20_0_ ( .in(spi_ss_in_bbank[0]),
     .out(spi_ss_in_bbankd[0]));
bram_bufferx16 I8_7_ ( .in(spi_ss_in_r[7]), .out(spi_ss_in_rd[7]));
bram_bufferx16 I8_6_ ( .in(spi_ss_in_r[6]), .out(spi_ss_in_rd[6]));
bram_bufferx16 I8_5_ ( .in(spi_ss_in_r[5]), .out(spi_ss_in_rd[5]));
bram_bufferx16 I8_4_ ( .in(spi_ss_in_r[4]), .out(spi_ss_in_rd[4]));
bram_bufferx16 I8_3_ ( .in(spi_ss_in_r[3]), .out(spi_ss_in_rd[3]));
bram_bufferx16 I8_2_ ( .in(spi_ss_in_r[2]), .out(spi_ss_in_rd[2]));
bram_bufferx16 I8_1_ ( .in(spi_ss_in_r[1]), .out(spi_ss_in_rd[1]));
ml_cram_logic Iml_cram_logic ( .smc_wwlwrt_en(net246),
     .smc_wset_precgnd(net248), .smc_write(smc_write),
     .cram_pgateoff(cram_pgateoff), .smc_wcram_rst(net252),
     .smc_rwl_en(net254), .smc_rrst_pullwlen(net256),
     .smc_rpull_b(net257), .smc_rprec(net258), .smc_read(net260),
     .smc_clk(net290), .por(core_por_bb), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_rst(cram_rst),
     .cram_pullup_b(cram_pullup_b), .cram_prec(cram_prec),
     .cram_vddoff(cram_vddoff), .smc_seq_rst(net253),
     .smc_clk_out(smc_clk_out), .smc_wwlwrt_dis(net247),
     .smc_wset_prec(net249));

endmodule
// Library - NVCM, Cell - ml_lshv_6v_hold, View - schematic
// LAST TIME SAVED: Dec 20 11:32:52 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_lshv_6v_hold ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M7 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(GND_), .G(vddp_tieh), .S(net132));
nch_25  M15 ( .D(net132), .B(GND_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(GND_), .G(vddp_tieh), .S(net140));
nch_25  M14 ( .D(net140), .B(GND_), .G(sel_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hv_inv, View - schematic
// LAST TIME SAVED: Jan 21 18:15:24 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_hv_inv ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
pch_25  M39 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM, Cell - ml_hv_ls_inv, View - schematic
// LAST TIME SAVED: Jan  8 14:11:13 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_hv_ls_inv ( in_hv, out_b_hv, sel_25, sel_b_25, vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_lshv_6v_hold Ishv_6v_hold ( .vddp_tieh(vddp_tieh), .out_b_hv(net61),
     .in_hv(in_hv), .sel_b_25(sel_b_25), .sel_25(sel_25),
     .out_hv(sel_hv));
ml_hv_inv Ihv_inv ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));

endmodule
// Library - tsmcN65lo, Cell - nand3_25, View - schematic
// LAST TIME SAVED: Mar 29 20:19:50 2006
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module nand3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(net21), .B(Gb), .G(C), .S(G));
nch_25  M2 ( .D(net25), .B(Gb), .G(B), .S(net21));
nch_25  NM1 ( .D(Y), .B(Gb), .G(A), .S(net25));
pch_25  PM1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M1 ( .D(Y), .B(Pb), .G(C), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(P));

endmodule
// Library - io, Cell - PVDD2POC, View - schematic
// LAST TIME SAVED: Jul 28 17:15:17 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module PVDD2POC ( VDDPST );
input  VDDPST;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - tsmcN65lo, Cell - nor3_25, View - schematic
// LAST TIME SAVED: Mar 29 20:26:16 2006
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module nor3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M2 ( .D(Y), .B(Gb), .G(A), .S(G));
nch_25  M3 ( .D(Y), .B(Gb), .G(C), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(B), .S(G));
pch_25  M1 ( .D(Y), .B(Pb), .G(C), .S(net16));
pch_25  PM1 ( .D(net12), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(net16), .B(Pb), .G(B), .S(net12));

endmodule
// Library - NVCM, Cell - ml_ls_vdd2vdd25, View - schematic
// LAST TIME SAVED: Apr  4 14:26:57 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
pch_25  M13 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
pch_25  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));
pch_25  M6 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
nch_25  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
nch_25  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));

endmodule
// Library - tsmcN65lo, Cell - inv_25, View - schematic
// LAST TIME SAVED: Mar 29 20:14:12 2006
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module inv_25 ( OUT, G, Gb, IN, P, Pb );
output  OUT;

input  G, Gb, IN, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  NM1 ( .D(OUT), .B(Gb), .G(IN), .S(G));
pch_25  PM1 ( .D(OUT), .B(Pb), .G(IN), .S(P));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tielow, View - schematic
// LAST TIME SAVED: May  8 16:23:59 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module vdd_tielow ( gnd_tiel );
inout  gnd_tiel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(gnd_tiel), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(net9), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_chip_spare, View - schematic
// LAST TIME SAVED: Sep 11 18:02:11 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_chip_spare (  );supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(net96), .B(net85), .G(net286), .S(net85));
pch_25  M5 ( .D(net85), .B(net123), .G(net114), .S(net123));
pch_25  M3 ( .D(net108), .B(net89), .G(net316), .S(net89));
pch_25  M2 ( .D(net89), .B(net126), .G(net119), .S(net126));
nch_25  M7 ( .D(net100), .B(GND_), .G(net286), .S(gnd_));
nch_25  M1 ( .D(net96), .B(GND_), .G(net121), .S(net100));
nch_25  M6 ( .D(net104), .B(GND_), .G(net316), .S(gnd_));
nch_25  M4 ( .D(net108), .B(GND_), .G(net121), .S(net104));
ml_hv_ls_inv I132 ( .sel_b_25(net316), .sel_25(net405),
     .out_b_hv(net119), .in_hv(net126), .vddp_tieh(net121));
ml_hv_ls_inv Iml_hv_ls_inv_vppt ( .sel_b_25(net286), .sel_25(net404),
     .out_b_hv(net114), .in_hv(net123), .vddp_tieh(net121));
rppolywo_m  R8 ( .MINUS(vddp_), .PLUS(net123), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(vddp_), .PLUS(net126), .BULK(gnd_));
nand3_25 I257 ( .B(net0373), .A(net0373), .Y(net0397), .C(net0373),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I256 ( .B(net0381), .A(net0381), .Y(net0373), .C(net0381),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I255 ( .B(net215), .A(net215), .Y(net0381), .C(net215),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I248 ( .B(net0397), .A(net0397), .Y(net0405), .C(net0397),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I247 ( .B(net0405), .A(net0405), .Y(net0413), .C(net0405),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I245 ( .B(net0413), .A(net0413), .Y(net0421), .C(net0413),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I244 ( .B(net0421), .A(net0421), .Y(net0453), .C(net0421),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I231 ( .B(net0453), .A(net0453), .Y(net0445), .C(net0453),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I233 ( .B(net0437), .A(net0437), .Y(net0429), .C(net0437),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I234 ( .B(net0429), .A(net0429), .Y(net0595), .C(net0429),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I232 ( .B(net0445), .A(net0445), .Y(net0437), .C(net0445),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nor3_25 I215 ( .B(net0460), .A(net0460), .C(net0460), .Y(net0594),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I214 ( .B(net0468), .A(net0468), .C(net0468), .Y(net0460),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I212 ( .B(net0476), .A(net0476), .C(net0476), .Y(net0468),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I211 ( .B(net160), .A(net160), .C(net160), .Y(net0492),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I209 ( .B(net0500), .A(net0500), .C(net0500), .Y(net0476),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I42 ( .B(net191), .A(net191), .C(net191), .Y(net160), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I78 ( .B(net199), .A(net199), .C(net199), .Y(net191), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I83 ( .B(net207), .A(net207), .C(net207), .Y(net199), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I84 ( .B(net215), .A(net215), .C(net215), .Y(net207), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I210 ( .B(net0492), .A(net0492), .C(net0492), .Y(net0500),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
inv_hvt I120 ( .A(net253), .Y(net249));
inv_hvt I119 ( .A(net231), .Y(net253));
inv_hvt I118 ( .A(net231), .Y(net258));
inv_hvt I117 ( .A(net258), .Y(net254));
inv_hvt I319 ( .A(net263), .Y(net259));
inv_hvt I323 ( .A(net231), .Y(net263));
inv_hvt I57 ( .A(net231), .Y(net268));
inv_hvt I58 ( .A(net268), .Y(net264));
ml_ls_vdd2vdd25 I122 ( .in(net249), .sup(vddp_), .out_vddio_b(net291),
     .out_vddio(net252), .in_b(net253));
ml_ls_vdd2vdd25 I121 ( .in(net254), .sup(vddp_), .out_vddio_b(net297),
     .out_vddio(net257), .in_b(net258));
ml_ls_vdd2vdd25 I335 ( .in(net259), .sup(vddp_), .out_vddio_b(net303),
     .out_vddio(net262), .in_b(net263));
ml_ls_vdd2vdd25 I56 ( .in(net264), .sup(vddp_), .out_vddio_b(net309),
     .out_vddio(net267), .in_b(net268));
inv_25 I126 ( .IN(net291), .OUT(net271), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I125 ( .IN(net297), .OUT(net272), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I139 ( .IN(net405), .OUT(net316), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(net404), .OUT(net286), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I384 ( .IN(net303), .OUT(net274), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I54 ( .IN(net309), .OUT(net273), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nand3_hvt I185 ( .Y(net0665), .B(net0661), .C(net0661), .A(net0661));
nand3_hvt I186 ( .Y(net0661), .B(net0657), .C(net0657), .A(net0657));
nand3_hvt I187 ( .Y(net0657), .B(net0653), .C(net0653), .A(net0653));
nand3_hvt I188 ( .Y(net0653), .B(net0649), .C(net0649), .A(net0649));
nand3_hvt I183 ( .Y(net0649), .B(net281), .C(net281), .A(net281));
nand3_hvt I246 ( .Y(net328), .B(net324), .C(net324), .A(net324));
nand3_hvt I61 ( .Y(net332), .B(net328), .C(net328), .A(net328));
nand3_hvt I62 ( .Y(net336), .B(net332), .C(net332), .A(net332));
nand3_hvt I63 ( .Y(net340), .B(net336), .C(net336), .A(net336));
nand3_hvt I64 ( .Y(net360), .B(net340), .C(net340), .A(net340));
nand3_hvt I104 ( .Y(net281), .B(net344), .C(net344), .A(net344));
nand3_hvt I105 ( .Y(net344), .B(net348), .C(net348), .A(net348));
nand3_hvt I106 ( .Y(net348), .B(net352), .C(net352), .A(net352));
nand3_hvt I107 ( .Y(net352), .B(net356), .C(net356), .A(net356));
nand3_hvt I108 ( .Y(net356), .B(net360), .C(net360), .A(net360));
nand3_hvt I184 ( .Y(net0596), .B(net0665), .C(net0665), .A(net0665));
nor3_hvt I177 ( .B(net0732), .Y(net0728), .A(net0732), .C(net0732));
nor3_hvt I178 ( .B(net0728), .Y(net0724), .A(net0728), .C(net0728));
nor3_hvt I179 ( .B(net0724), .Y(net0720), .A(net0724), .C(net0724));
nor3_hvt I180 ( .B(net0720), .Y(net0716), .A(net0720), .C(net0720));
nor3_hvt I181 ( .B(net0716), .Y(net0712), .A(net0716), .C(net0716));
nor3_hvt I182 ( .B(net0712), .Y(net0597), .A(net0712), .C(net0712));
nor3_hvt I65 ( .B(net363), .Y(net383), .A(net363), .C(net363));
nor3_hvt I70 ( .B(net367), .Y(net363), .A(net367), .C(net367));
nor3_hvt I71 ( .B(net371), .Y(net367), .A(net371), .C(net371));
nor3_hvt I72 ( .B(net375), .Y(net371), .A(net375), .C(net375));
nor3_hvt I73 ( .B(net379), .Y(net375), .A(net379), .C(net379));
nor3_hvt I99 ( .B(net383), .Y(net387), .A(net383), .C(net383));
nor3_hvt I100 ( .B(net387), .Y(net391), .A(net387), .C(net387));
nor3_hvt I101 ( .B(net391), .Y(net395), .A(net391), .C(net391));
nor3_hvt I102 ( .B(net395), .Y(net399), .A(net395), .C(net395));
nor3_hvt I103 ( .B(net399), .Y(net0732), .A(net399), .C(net399));
vddp_tiehigh I140 ( .vddp_tieh(net121));
vdd_tielow I154 ( .gnd_tiel(net405));
vdd_tielow I155 ( .gnd_tiel(net404));
vdd_tielow I153 ( .gnd_tiel(net231));
vdd_tielow I146 ( .gnd_tiel(net215));
vdd_tielow I145 ( .gnd_tiel(net324));
vdd_tielow I144 ( .gnd_tiel(net379));

endmodule
// Library - tsmcN65lo, Cell - nand2_25, View - schematic
// LAST TIME SAVED: Mar 29 20:17:19 2006
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module nand2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(net16), .B(Gb), .G(B), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(A), .S(net16));
pch_25  M2 ( .D(Y), .B(Pb), .G(B), .S(P));
pch_25  PM1 ( .D(Y), .B(Pb), .G(A), .S(P));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr, View - schematic
// LAST TIME SAVED: Feb 25 14:20:48 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr ( wr, gwl_wr_25, s_25, wr_sup_25 );
output  wr;

input  gwl_wr_25, s_25, wr_sup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_25 I59 ( .A(gwl_wr_25), .Y(net27), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(s_25));
inv_25 I38 ( .IN(net27), .OUT(wr), .P(wr_sup_25), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr_x4, View - schematic
// LAST TIME SAVED: Jan 21 18:09:38 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x4 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  gwl_wr_25, wr_sup_25;

output [3:0]  wr;

input [3:0]  s_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr Iml_lwldrv_2 ( .gwl_wr_25(gwl_wr_25), .wr(wr[2]),
     .s_25(s_25[2]), .wr_sup_25(wr_sup_25));
ml_rock_lwldrv_wr Iml_lwldrv_1 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[1]), .wr(wr[1]));
ml_rock_lwldrv_wr Iml_lwldrv_3 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3]), .wr(wr[3]));
ml_rock_lwldrv_wr Iml_lwldrv_0 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[0]), .wr(wr[0]));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr_x27_1f, View - schematic
// LAST TIME SAVED: Jan 20 17:28:59 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x27_1f ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  wr_sup_25;

output [107:0]  wr;

input [26:0]  gwl_wr_25;
input [3:0]  s_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_26_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[107:104]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[26]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_25_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[103:100]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[25]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_24_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[99:96]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[24]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_23_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[95:92]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[23]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_22_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[91:88]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[22]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_21_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[87:84]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[21]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_20_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[83:80]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[20]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_19_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[79:76]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[19]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_18_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[75:72]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[18]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_17_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[71:68]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[17]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_16_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[67:64]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[16]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_15_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[63:60]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[15]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_14_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[59:56]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[14]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_13_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[55:52]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[13]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_12_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[51:48]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[12]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_11_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[47:44]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[11]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_10_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[43:40]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[10]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_9_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[39:36]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[9]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_8_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[35:32]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[8]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_7_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[31:28]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[7]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_6_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[27:24]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[6]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_5_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[23:20]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[5]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_4_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[19:16]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[4]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_3_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[15:12]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[3]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_2_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[11:8]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[2]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_1_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[7:4]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[1]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_0_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[3:0]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[0]));

endmodule
// Library - NVCM, Cell - ml_ls_vddp2vpxa, View - schematic
// LAST TIME SAVED: Dec 30 20:36:23 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_ls_vddp2vpxa ( out_33, out_b_33, sup, in_25, in_b_25 );
output  out_33, out_b_33;

inout  sup;

input  in_25, in_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(out_b_33), .B(sup), .G(in_25), .S(net29));
pch_25  M13 ( .D(out_33), .B(sup), .G(in_b_25), .S(net33));
pch_25  M4 ( .D(net29), .B(sup), .G(out_33), .S(sup));
pch_25  M6 ( .D(net33), .B(sup), .G(out_b_33), .S(sup));
nch_25  M9 ( .D(out_33), .B(gnd_), .G(in_b_25), .S(gnd_));
nch_25  M15 ( .D(out_b_33), .B(gnd_), .G(in_25), .S(gnd_));

endmodule
// Library - io, Cell - PVDD2DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:14:57 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module PVDD2DGZ ( VDDPST );
input  VDDPST;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - tsmcN65lo, Cell - nor2_25, View - schematic
// LAST TIME SAVED: Mar 29 20:24:25 2006
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module nor2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(Y), .B(Gb), .G(A), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(B), .S(G));
pch_25  PM1 ( .D(net15), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(net15));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_gwhv, View - schematic
// LAST TIME SAVED: May 16 11:27:16 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_rock_lwldrv_gwhv ( gwp_hv, gwp_sup_hv, gwl_25, gwl_25_b,
     vddp_tieh );
output  gwp_hv;

inout  gwp_sup_hv;

input  gwl_25, gwl_25_b, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M10 ( .D(net0129), .B(gnd_), .G(vddp_tieh), .S(net050));
nch_25  M12 ( .D(gwp_hv), .B(gnd_), .G(vddp_tieh), .S(net034));
nch_25  M11 ( .D(net034), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M13 ( .D(net050), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M14 ( .D(net054), .B(gnd_), .G(vddp_tieh), .S(net058));
nch_25  M15 ( .D(net058), .B(gnd_), .G(gwl_25), .S(gnd_));
pch_25  M6 ( .D(net067), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M16 ( .D(gwp_hv), .B(net067), .G(gwl_25_b), .S(net067));
pch_25  M5 ( .D(net054), .B(net087), .G(gwl_25), .S(net087));
pch_25  M8 ( .D(net087), .B(gwp_sup_hv), .G(net0129), .S(gwp_sup_hv));
pch_25  M9 ( .D(net091), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M7 ( .D(net0129), .B(net091), .G(gwl_25_b), .S(net091));

endmodule
// Library - NVCM, Cell - ml_gwl_drv, View - schematic
// LAST TIME SAVED: Apr 30 15:58:52 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_gwl_drv ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25,
     radd_1_25, radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );
output  gwl_b_25, gwl_wr_25, gwp_hv;

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25, radd_1_25,
     radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ls_vddp2vpxa I99 ( .in_25(gwlb_25), .sup(gwl_b_sup_25),
     .in_b_25(gwlb_b_25), .out_33(out_33), .out_b_33(net053));
nor3_25 I76 ( .C(net84), .A(net68), .Y(dec_sel_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(net76));
nor2_25 I111 ( .A(net096), .Y(gwlb_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_dis_25));
nor2_25 I79 ( .A(wr_dis_25), .Y(gwl_wr_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(net056));
nor2_25 I117 ( .A(dec_sel_25), .Y(net096), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_en_25));
nor2_25 I82 ( .A(dec_sel_25), .Y(net058), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_frcen_25));
nor2_25 I85 ( .A(net058), .Y(gwl_wp_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_dis_25));
nor2_25 I59 ( .B(dec_sel_25), .A(wr_frcen_25), .Y(net056), .P(vddp_),
     .Pb(vddp_), .Gb(gnd_), .G(gnd_));
ml_rock_lwldrv_gwhv Iml_rock_lwldrv_gwhv ( .gwp_sup_hv(gwp_sup_hv),
     .vddp_tieh(vddp_tieh), .gwp_hv(gwp_hv), .gwl_25(gwl_wp_25),
     .gwl_25_b(gwl_wp_b_25));
nand3_25 I44 ( .B(radd_4_25), .A(radd_5_25), .Y(net76), .C(radd_3_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I47 ( .B(radd_1_25), .A(radd_2_25), .Y(net84), .C(radd_0_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I104 ( .B(gwlgrpsel_25), .A(gwlgrpsel_25), .Y(net68),
     .C(radd_6_25), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
inv_25 I38 ( .IN(gwl_wp_25), .OUT(gwl_wp_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I100 ( .IN(out_33), .OUT(gwl_b_25), .P(gwl_b_sup_25),
     .Pb(gwl_b_sup_25), .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(gwlb_25), .OUT(gwlb_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_gwl_drv_x27_1f, View - schematic
// LAST TIME SAVED: Feb 11 11:36:23 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_gwl_drv_x27_1f ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25,
     gnv2_b_25, gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25,
     gnv5_b_25, gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1,
     gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25, gnv2_b_25,
     gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25, gnv5_b_25,
     gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1, gwl_misc_25,
     gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

output [26:0]  gwl_b_25;
output [26:0]  gwp_hv;
output [26:0]  gwl_wr_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_gwl_drv Igwl_drv_25_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[25]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[25]), .gwl_wr_25(gwl_wr_25[25]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_24_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[24]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[24]), .gwl_wr_25(gwl_wr_25[24]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_23_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[23]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[23]), .gwl_wr_25(gwl_wr_25[23]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_22_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[22]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[22]), .gwl_wr_25(gwl_wr_25[22]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_21_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[21]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[21]), .gwl_wr_25(gwl_wr_25[21]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_20_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[20]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[20]), .gwl_wr_25(gwl_wr_25[20]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_19_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[19]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[19]), .gwl_wr_25(gwl_wr_25[19]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_18_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[18]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[18]), .gwl_wr_25(gwl_wr_25[18]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_17_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[17]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[17]), .gwl_wr_25(gwl_wr_25[17]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_16_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[16]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[16]), .gwl_wr_25(gwl_wr_25[16]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_misc_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[26]),
     .radd_0_25(vddp_tieh), .radd_1_25(vddp_tieh),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_misc_25),
     .gwp_hv(gwp_hv[26]), .gwl_wr_25(gwl_wr_25[26]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_15_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[15]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[15]), .gwl_wr_25(gwl_wr_25[15]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_14_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[14]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[14]), .gwl_wr_25(gwl_wr_25[14]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_13_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[13]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[13]), .gwl_wr_25(gwl_wr_25[13]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_12_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[12]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[12]), .gwl_wr_25(gwl_wr_25[12]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_11_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[11]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[11]), .gwl_wr_25(gwl_wr_25[11]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_10_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[10]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[10]), .gwl_wr_25(gwl_wr_25[10]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_9_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[9]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[9]), .gwl_wr_25(gwl_wr_25[9]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_8_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[8]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[8]),
     .gwl_wr_25(gwl_wr_25[8]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_7_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[7]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[7]),
     .gwl_wr_25(gwl_wr_25[7]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_6_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[6]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[6]),
     .gwl_wr_25(gwl_wr_25[6]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_5_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[5]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[5]),
     .gwl_wr_25(gwl_wr_25[5]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_4_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[4]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[4]),
     .gwl_wr_25(gwl_wr_25[4]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_3_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[3]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[3]),
     .gwl_wr_25(gwl_wr_25[3]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_2_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[2]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[2]),
     .gwl_wr_25(gwl_wr_25[2]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_1_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[1]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[1]),
     .gwl_wr_25(gwl_wr_25[1]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[0]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_b_25),
     .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[0]), .gwl_wr_25(gwl_wr_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM, Cell - ml_gwlwr_1f, View - schematic
// LAST TIME SAVED: Jan 20 17:29:06 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_gwlwr_1f ( gwl_b_25, gwp_hv, wr, gwl_b_sup_25, gwp_sup_hv,
     gnv_25, gnv_b_25, gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25,
     gwl_red_25, gwlb_dis_25, gwlb_en_25, s_25, vddp_tieh, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, wr_sup_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wr_sup_25;

output [107:0]  wr;
output [26:0]  gwl_b_25;
output [26:0]  gwp_hv;

input [3:0]  s_25;
input [1:0]  gred_25;
input [5:0]  gnv_b_25;
input [1:0]  gred_b_25;
input [5:0]  gnv_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [26:0]  gwl_wr_25;



ml_rock_lwldrv_wr_x27_1f Iml_rock_lwldrv_wr_x27_1f (
     .gwl_wr_25(gwl_wr_25[26:0]), .wr(wr[107:0]),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3:0]));
ml_gwl_drv_x27_1f Iml_gwl_drv_x27_1f ( .gwp_hv(gwp_hv[26:0]),
     .gwl_wr_25(gwl_wr_25[26:0]), .gwl_b_25(gwl_b_25[26:0]),
     .gwlb_en_25(gwlb_en_25), .gwlb_dis_25(gwlb_dis_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25_1(gred_b_25[1]), .gred_b_25_0(gred_b_25[0]),
     .gred_25_1(gred_25[1]), .gred_25_0(gred_25[0]),
     .gnv5_b_25(gnv_b_25[5]), .gnv5_25(gnv_25[5]),
     .gnv4_b_25(gnv_b_25[4]), .gnv4_25(gnv_25[4]),
     .gnv3_b_25(gnv_b_25[3]), .gnv3_25(gnv_25[3]),
     .gnv2_b_25(gnv_b_25[2]), .gnv2_25(gnv_25[2]),
     .gnv1_b_25(gnv_b_25[1]), .gnv1_25(gnv_25[1]),
     .gnv0_b_25(gnv_b_25[0]), .gnv0_25(gnv_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));

endmodule
// Library - NVCM, Cell - ml_hv_invx3_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:19:36 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_hv_invx3_enhance ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh
     );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM, Cell - ml_lshv_6v_switch_enhance, View - schematic
// LAST TIME SAVED: Apr 30 14:46:53 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_lshv_6v_switch_enhance ( out_b_hv, out_hv, in_hv, sel_25,
     sel_b_25, vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
nch_25  M11 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hv_ls_inv_hotsw_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:16:13 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw_enhance ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3_enhance Ihv_invx3 ( .vddp_tieh(vddp_tieh),
     .out_b_hv(out_b_hv), .sel_25(sel_25), .in_hv(in_hv),
     .sel_hv(sel_hv));
ml_lshv_6v_switch_enhance Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM, Cell - ml_hv_hotswitch_enhance, View - schematic
// LAST TIME SAVED: Jan 23 14:29:21 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_hv_hotswitch_enhance ( hv_in_hv, hv_out_hv, selhv_25,
     vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));
nch_25  M7 ( .D(net12), .B(GND_), .G(selhv_25), .S(net15));
nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
nch_25  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
pch_25  M0 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_hotswitch_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:28:27 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch_enhance ( hvin_a_hv, hvin_b_hv, out_hv,
     sel_hv_a_25, sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch_enhance Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - io, Cell - lefbank_1k_july16, View - schematic
// LAST TIME SAVED: Jul 16 11:35:48 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module lefbank_1k_july16 ( in, pad, oen, out, ren );



output [25:0]  in;

inout [25:0]  pad;

input [25:0]  oen;
input [25:0]  out;
input [25:0]  ren;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



PDUW08DGZ I63_7_ ( .PAD(pad[7]), .C(in[7]), .OEN(oen[7]), .I(out[7]),
     .REN(ren[7]));
PDUW08DGZ I63_6_ ( .PAD(pad[6]), .C(in[6]), .OEN(oen[6]), .I(out[6]),
     .REN(ren[6]));
PDUW08DGZ I61_5_ ( .PAD(pad[5]), .C(in[5]), .OEN(oen[5]), .I(out[5]),
     .REN(ren[5]));
PDUW08DGZ I61_4_ ( .PAD(pad[4]), .C(in[4]), .OEN(oen[4]), .I(out[4]),
     .REN(ren[4]));
PDUW08DGZ I61_3_ ( .PAD(pad[3]), .C(in[3]), .OEN(oen[3]), .I(out[3]),
     .REN(ren[3]));
PDUW08DGZ I61_2_ ( .PAD(pad[2]), .C(in[2]), .OEN(oen[2]), .I(out[2]),
     .REN(ren[2]));
PDUW08DGZ I61_1_ ( .PAD(pad[1]), .C(in[1]), .OEN(oen[1]), .I(out[1]),
     .REN(ren[1]));
PDUW08DGZ I61_0_ ( .PAD(pad[0]), .C(in[0]), .OEN(oen[0]), .I(out[0]),
     .REN(ren[0]));
PDUW08DGZ I92_21_ ( .PAD(pad[21]), .C(in[21]), .OEN(oen[21]),
     .I(out[21]), .REN(ren[21]));
PDUW08DGZ I92_20_ ( .PAD(pad[20]), .C(in[20]), .OEN(oen[20]),
     .I(out[20]), .REN(ren[20]));
PDUW08DGZ I92_19_ ( .PAD(pad[19]), .C(in[19]), .OEN(oen[19]),
     .I(out[19]), .REN(ren[19]));
PDUW08DGZ I92_18_ ( .PAD(pad[18]), .C(in[18]), .OEN(oen[18]),
     .I(out[18]), .REN(ren[18]));
PDUW08DGZ I92_17_ ( .PAD(pad[17]), .C(in[17]), .OEN(oen[17]),
     .I(out[17]), .REN(ren[17]));
PDUW08DGZ I92_16_ ( .PAD(pad[16]), .C(in[16]), .OEN(oen[16]),
     .I(out[16]), .REN(ren[16]));
PDUW08DGZ I102_11_ ( .PAD(pad[11]), .C(in[11]), .OEN(oen[11]),
     .I(out[11]), .REN(ren[11]));
PDUW08DGZ I102_10_ ( .PAD(pad[10]), .C(in[10]), .OEN(oen[10]),
     .I(out[10]), .REN(ren[10]));
PDUW08DGZ I102_9_ ( .PAD(pad[9]), .C(in[9]), .OEN(oen[9]), .I(out[9]),
     .REN(ren[9]));
PDUW08DGZ I102_8_ ( .PAD(pad[8]), .C(in[8]), .OEN(oen[8]), .I(out[8]),
     .REN(ren[8]));
PDUW08DGZ I101_15_ ( .PAD(pad[15]), .C(in[15]), .OEN(oen[15]),
     .I(out[15]), .REN(ren[15]));
PDUW08DGZ I101_14_ ( .PAD(pad[14]), .C(in[14]), .OEN(oen[14]),
     .I(out[14]), .REN(ren[14]));
PDUW08DGZ I60_25_ ( .PAD(pad[25]), .C(in[25]), .OEN(oen[25]),
     .I(out[25]), .REN(ren[25]));
PDUW08DGZ I60_24_ ( .PAD(pad[24]), .C(in[24]), .OEN(oen[24]),
     .I(out[24]), .REN(ren[24]));
PDUW08DGZ I60_23_ ( .PAD(pad[23]), .C(in[23]), .OEN(oen[23]),
     .I(out[23]), .REN(ren[23]));
PDUW08DGZ I60_22_ ( .PAD(pad[22]), .C(in[22]), .OEN(oen[22]),
     .I(out[22]), .REN(ren[22]));
PDUW08DGZ I58_13_ ( .PAD(pad[13]), .C(in[13]), .OEN(oen[13]),
     .I(out[13]), .REN(ren[13]));
PDUW08DGZ I58_12_ ( .PAD(pad[12]), .C(in[12]), .OEN(oen[12]),
     .I(out[12]), .REN(ren[12]));
PVSS3DGZ I98 ( .VSS(gnd_));
PVSS3DGZ I85_1_ ( .VSS(gnd_));
PVSS3DGZ I85_0_ ( .VSS(gnd_));
PVSS3DGZ I97_1_ ( .VSS(gnd_));
PVSS3DGZ I97_0_ ( .VSS(gnd_));
PVSS3DGZ I90_1_ ( .VSS(gnd_));
PVSS3DGZ I90_0_ ( .VSS(gnd_));
PVSS3DGZ I100_1_ ( .VSS(gnd_));
PVSS3DGZ I100_0_ ( .VSS(gnd_));
PVDD1DGZ I87_1_ ( .VDD(vdd_));
PVDD1DGZ I87_0_ ( .VDD(vdd_));
PVDD1DGZ I99 ( .VDD(vdd_));
PVDD2POC I93 ( .VDDPST(vddio_leftbank));
PVDD2DGZ I91_1_ ( .VDDPST(vddio_leftbank));
PVDD2DGZ I91_0_ ( .VDDPST(vddio_leftbank));
PVDD2DGZ I95_1_ ( .VDDPST(vddio_leftbank));
PVDD2DGZ I95_0_ ( .VDDPST(vddio_leftbank));
PVDD2DGZ I94 ( .VDDPST(vddio_leftbank));

endmodule
// Library - sbtlibn65lp, Cell - oai22x2_hvt, View - schematic
// LAST TIME SAVED: Jan 24 13:53:38 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module oai22x2_hvt ( Y, A0, A1, B0, B1 );
output  Y;

input  A0, A1, B0, B1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(Y), .B(GND_), .G(A0), .S(net024));
nch_hvt  M8 ( .D(Y), .B(GND_), .G(A1), .S(net024));
nch_hvt  M10 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
pch_hvt  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M4 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
pch_hvt  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_pump_a_clkdly, View - schematic
// LAST TIME SAVED: Feb 11 09:24:13 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module ml_pump_a_clkdly ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(net66), .S(vdd_));
pch_hvt  M0 ( .D(vdd_), .B(vdd_), .G(net62), .S(vdd_));
inv_hvt I206 ( .A(in), .Y(net66));
inv_hvt I204 ( .A(net64), .Y(net62));
inv_hvt I205 ( .A(net66), .Y(net64));
inv_hvt I207 ( .A(net70), .Y(out));
inv_hvt I208 ( .A(net62), .Y(net70));

endmodule
// Library - sbtlibn65lp, Cell - anor31_hvt, View - schematic
// LAST TIME SAVED: Feb 13 14:15:10 2008
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module anor31_hvt ( Y, A, B, C, D );
output  Y;

input  A, B, C, D;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(Y), .B(gnd_), .G(A), .S(net23));
nch_hvt  M8 ( .D(net030), .B(gnd_), .G(C), .S(gnd_));
nch_hvt  M6 ( .D(net23), .B(gnd_), .G(B), .S(net030));
nch_hvt  M7 ( .D(Y), .B(gnd_), .G(D), .S(gnd_));
pch_hvt  M5 ( .D(Y), .B(vdd_), .G(D), .S(net35));
pch_hvt  M4 ( .D(net35), .B(vdd_), .G(A), .S(vdd_));
pch_hvt  M3 ( .D(net35), .B(vdd_), .G(B), .S(vdd_));
pch_hvt  M2 ( .D(net35), .B(vdd_), .G(C), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_logic, View - schematic
// LAST TIME SAVED: Mar  4 15:44:43 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_logic ( gnv, gred, gwl_misc, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, s, sa_trim, saen, testdec_en_b, testdec_even_b,
     testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd, fsm_coladd, fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_trow, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_dma, tm_testdec, tm_testdec_wr );
output  gwl_misc, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, saen, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [5:0]  gnv;
output [1:0]  gred;
output [3:0]  s;
output [2:0]  sa_trim;

input [7:0]  fsm_rowadd;
input [0:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_b;

wire  [5:0]  gnv_b;

wire  [2:0]  sa_trim_b;

wire  [1:0]  xadd_b;

wire  [1:0]  gred_b;

wire  [1:0]  xadd;

wire  [0:2]  net390;

wire  [0:1]  net386;



vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
anor21_hvt I109_1_ ( .A(net386[0]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I109_0_ ( .A(net386[1]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
oai22x2_hvt I93 ( .A1(fsm_rd), .Y(net196), .A0(fsm_pgmvfy),
     .B0(gnd_tiel), .B1(gnd_tiel));
ml_pump_a_clkdly I230 ( .in(net0231), .out(net0232));
ml_pump_a_clkdly I208 ( .in(net200), .out(net201));
ml_pump_a_clkdly I202 ( .in(net202), .out(net203));
ml_pump_a_clkdly I198 ( .in(net204), .out(net205));
ml_pump_a_clkdly I207 ( .in(net206), .out(net207));
nor4_hvt I175 ( .D(fsm_tm_allwl_h), .B(fsm_pgmvfy), .Y(net211),
     .A(fsm_pgmvfy), .C(fsm_rd));
nor4_hvt I176 ( .D(testdec_wp), .B(fsm_nvcmen_b), .Y(net216),
     .A(fsm_wren_b), .C(net331));
nor4_hvt I218 ( .D(net282), .B(fsm_tm_allbl_l), .Y(net0258),
     .A(fsm_tm_allbl_l), .C(fsm_nvcmen_b));
nor4_hvt I191 ( .B(pgm_hvpulse), .Y(wrsup_2vdd_int), .D(fsm_nvcmen_b),
     .A(pgm_hvpulse), .C(testdec_wr));
nor4_hvt I171 ( .D(fsm_wpen_b), .B(fsm_nvcmen_b), .Y(net226),
     .A(testdec_wr), .C(fsm_tm_allwl_l));
nor2_hvt I233 ( .A(fsm_pgm), .B(fsm_pgmvfy), .Y(net0176));
nor2_hvt I228 ( .A(fsm_pgmdisc), .B(fsm_pgmhv), .Y(net0231));
nor2_hvt I231 ( .A(net0258), .B(tm_testdec), .Y(pgminhi_dmmy_b));
nor2_hvt I165 ( .B(fsm_nv_sisi_ui), .Y(x1_desel_b),
     .A(fsm_nv_rri_trim));
nor2_hvt I131 ( .B(tm_testdec_wr), .A(testdec_en_b), .Y(testdec_en));
nor2_hvt I186 ( .A(fsm_pgmvfy), .B(fsm_pgm_b), .Y(stress2));
nor2_hvt I216 ( .A(fsm_nvcmen_b), .B(tm_dma), .Y(saen));
nor2_hvt I203 ( .A(net203), .B(net351), .Y(gwlbsup_vpxa));
nor2_hvt I209 ( .A(net207), .B(net246), .Y(gwphv_vppint));
nor2_hvt I214 ( .A(net0232), .B(fsm_nvcmen_b), .Y(net246));
nor2_hvt I210 ( .A(net359), .B(net201), .Y(gwphv_vddp));
nor2_hvt I226 ( .A(net0288), .B(net0390), .Y(gwlb_en));
nor2_hvt I201 ( .A(net196), .B(net205), .Y(gwlbsup_vddp));
nor3_hvt I182 ( .B(fsm_tm_allwl_l), .Y(net330), .A(fsm_tm_allwl_l),
     .C(fsm_tm_allwl_l));
nor3_hvt I105 ( .B(fsm_tm_allwl_h), .Y(net0288), .A(fsm_tm_allwl_h),
     .C(fsm_tm_allwl_h));
nor3_hvt I162 ( .Y(net0274), .B(fsm_tm_trow), .C(fsm_nv_sisi_ui),
     .A(fsm_nv_rri_trim));
anor31_hvt I121_3_ ( .A(net365), .D(net345), .B(xadd[1]), .Y(s_b[3]),
     .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net365), .D(net345), .B(xadd[1]), .Y(s_b[2]),
     .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net365), .D(net345), .B(xadd_b[1]), .Y(s_b[1]),
     .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net365), .D(net345), .B(xadd_b[1]), .Y(s_b[0]),
     .C(xadd_b[0]));
nand3_hvt I167 ( .B(fsm_nvcmen), .Y(gwlb_dis), .A(net0332),
     .C(testwr_wpgnd_b));
nand3_hvt I184 ( .Y(net274), .B(fsm_tm_allwl_h), .C(fsm_tm_allwl_h),
     .A(stress2));
nand3_hvt I125 ( .C(fsm_ymuxdis), .A(tm_testdec), .Y(testdec_prec_b),
     .B(fsm_rd));
nand3_hvt I195 ( .Y(net282), .B(net341), .C(fsm_lshven), .A(fsm_pgm));
nand3_hvt I154 ( .Y(net286), .B(fsm_pgm), .C(fsm_tm_allwl_h),
     .A(fsm_wren));
nand3_hvt I122 ( .A(fsm_nvcmen), .C(net307), .Y(net292),
     .B(tm_allwl_l_b));
nand2_hvt I170 ( .A(tm_testdec_wr), .Y(testwr_wpgnd_b),
     .B(tm_testdec));
nand2_hvt I188 ( .A(testdec_en), .Y(testdec_odd_b), .B(fsm_coladd[0]));
nand2_hvt I189 ( .A(net355), .Y(testdec_even_b), .B(testdec_en));
nand2_hvt I155 ( .A(net377), .Y(net307), .B(tm_testdec));
nand2_hvt I89 ( .A(fsm_rd), .Y(testdec_en_b), .B(tm_testdec));
inv_hvt I232 ( .A(net0176), .Y(net0365));
inv_hvt I174 ( .A(net211), .Y(wp_frcen));
inv_hvt I163 ( .A(net0274), .Y(gwl_misc));
inv_hvt I187 ( .A(fsm_pgm), .Y(fsm_pgm_b));
inv_hvt I178 ( .A(net307), .Y(testdec_wp));
inv_hvt I196 ( .A(net282), .Y(pgm_hvpulse));
inv_hvt I185 ( .A(net274), .Y(wr_frcen));
inv_hvt I206 ( .A(gwlbsup_vpxa), .Y(net204));
inv_hvt I177 ( .A(net216), .Y(wr_dis));
inv_hvt I183 ( .A(net330), .Y(net331));
inv_hvt I192 ( .A(wrsup_2vdd_int), .Y(net333));
inv_hvt I179 ( .A(fsm_wpen), .Y(fsm_wpen_b));
inv_hvt I194 ( .A(testwr_wpgnd_b), .Y(testdec_wr));
inv_hvt I212 ( .A(gwphv_vddp), .Y(net206));
inv_hvt I197 ( .A(fsm_pgmvfy), .Y(net341));
inv_hvt I205 ( .A(gwlbsup_vddp), .Y(net202));
inv_hvt I152 ( .A(net286), .Y(net345));
inv_hvt I120_5_ ( .A(gnv_b[5]), .Y(gnv[5]));
inv_hvt I120_4_ ( .A(gnv_b[4]), .Y(gnv[4]));
inv_hvt I120_3_ ( .A(gnv_b[3]), .Y(gnv[3]));
inv_hvt I120_2_ ( .A(gnv_b[2]), .Y(gnv[2]));
inv_hvt I120_1_ ( .A(gnv_b[1]), .Y(gnv[1]));
inv_hvt I120_0_ ( .A(gnv_b[0]), .Y(gnv[0]));
inv_hvt I172 ( .A(net226), .Y(wp_dis));
inv_hvt I204 ( .A(net196), .Y(net351));
inv_hvt I160_1_ ( .A(gred_b[1]), .Y(gred[1]));
inv_hvt I160_0_ ( .A(gred_b[0]), .Y(gred[0]));
inv_hvt I190 ( .A(fsm_coladd[0]), .Y(net355));
inv_hvt I150_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I150_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I215 ( .A(net246), .Y(net359));
inv_hvt I225 ( .A(pgm_hvpulse), .Y(net0390));
inv_hvt I213 ( .A(gwphv_vppint), .Y(net200));
inv_hvt I161_1_ ( .A(fsm_rowadd[3]), .Y(gred_b[1]));
inv_hvt I161_0_ ( .A(fsm_rowadd[2]), .Y(gred_b[0]));
inv_hvt I151 ( .A(net292), .Y(net365));
inv_hvt I119_5_ ( .A(fsm_rowadd[7]), .Y(gnv_b[5]));
inv_hvt I119_4_ ( .A(fsm_rowadd[6]), .Y(gnv_b[4]));
inv_hvt I119_3_ ( .A(fsm_rowadd[5]), .Y(gnv_b[3]));
inv_hvt I119_2_ ( .A(fsm_rowadd[4]), .Y(gnv_b[2]));
inv_hvt I119_1_ ( .A(fsm_rowadd[3]), .Y(gnv_b[1]));
inv_hvt I119_0_ ( .A(fsm_rowadd[2]), .Y(gnv_b[0]));
inv_hvt I157 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I153 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I193 ( .A(net333), .Y(wrsup_2vdd));
inv_hvt I181 ( .A(fsm_wren), .Y(fsm_wren_b));
inv_hvt I156 ( .A(tm_testdec_wr), .Y(net377));
inv_hvt I147_3_ ( .A(s_b[3]), .Y(s[3]));
inv_hvt I147_2_ ( .A(s_b[2]), .Y(s[2]));
inv_hvt I147_1_ ( .A(s_b[1]), .Y(s[1]));
inv_hvt I147_0_ ( .A(s_b[0]), .Y(s[0]));
inv_hvt I25_2_ ( .A(sa_trim_b[2]), .Y(sa_trim[2]));
inv_hvt I25_1_ ( .A(sa_trim_b[1]), .Y(sa_trim[1]));
inv_hvt I25_0_ ( .A(sa_trim_b[0]), .Y(sa_trim[0]));
inv_hvt I24_2_ ( .A(net390[0]), .Y(sa_trim_b[2]));
inv_hvt I24_1_ ( .A(net390[1]), .Y(sa_trim_b[1]));
inv_hvt I24_0_ ( .A(net390[2]), .Y(sa_trim_b[0]));
mux2_hvt I180_1_ ( .in1(fsm_rowadd[1]), .in0(fsm_rowadd[1]),
     .out(net386[0]), .sel(fsm_nv_rrow));
mux2_hvt I180_0_ ( .in1(fsm_rowadd[0]), .in0(fsm_rowadd[0]),
     .out(net386[1]), .sel(fsm_nv_rrow));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net390[0]), .sel(net0365));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net390[1]), .sel(net0365));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net390[2]), .sel(net0365));
mux2_hvt I221 ( .in1(fsm_wpen), .in0(fsm_wgnden), .out(net0332),
     .sel(pgm_hvpulse));

endmodule
// Library - NVCM, Cell - ml_hv_invx3, View - schematic
// LAST TIME SAVED: Jan 25 09:27:09 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_hv_invx3 ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM, Cell - ml_lshv_6v_switch, View - schematic
// LAST TIME SAVED: Feb  1 16:53:01 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_lshv_6v_switch ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
nch_25  M11 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hv_ls_inv_hotsw, View - schematic
// LAST TIME SAVED: Jan 24 11:18:40 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3 Ihv_invx3 ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));
ml_lshv_6v_switch Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM, Cell - ml_hv_hotswitch, View - schematic
// LAST TIME SAVED: Jan 25 09:27:57 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_hv_hotswitch ( hv_in_hv, hv_out_hv, selhv_25, vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));
nch_25  M7 ( .D(net12), .B(GND_), .G(selhv_25), .S(net15));
nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
nch_25  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
pch_25  M0 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_hotswitch, View - schematic
// LAST TIME SAVED: Jan 26 19:35:53 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch ( hvin_a_hv, hvin_b_hv, out_hv, sel_hv_a_25,
     sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - NVCM, Cell - ml_gwlwr_bldrv, View - schematic
// LAST TIME SAVED: Apr  9 11:04:12 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_gwlwr_bldrv ( bgr, bl_pgm_glb, bl_frc_gnd, fsm_din, fsm_pgm,
     fsm_pgmien, fsm_trim_ipp, tm_dma );
inout  bgr, bl_pgm_glb;

input  bl_frc_gnd, fsm_din, fsm_pgm, fsm_pgmien, tm_dma;

input [3:0]  fsm_trim_ipp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net0152;

wire  [0:3]  net0172;

wire  [0:3]  net0156;

wire  [0:7]  net0115;

wire  [0:1]  net0180;

wire  [0:1]  net0160;



nand2_hvt I71 ( .B(fsm_din), .A(fsm_pgmien), .Y(fsm_pgmien_b_buf));
nor2_hvt I121 ( .A(net086), .B(fsm_pgmien_b_buf), .Y(pgm_trim0_en));
nor2_hvt I114 ( .B(tm_dma), .Y(net0116), .A(tm_dma));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
nor4_hvt I105 ( .D(fsm_trim_ipp[0]), .B(fsm_trim_ipp[2]), .Y(net086),
     .A(fsm_trim_ipp[3]), .C(fsm_trim_ipp[1]));
nch_hvt  M36 ( .D(net0173), .B(GND_), .G(pgm_trim0_en), .S(net0107));
nch_hvt  M37 ( .D(net0107), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M31_7_ ( .D(net0115[0]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[0]));
nch_hvt  M31_6_ ( .D(net0115[1]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[1]));
nch_hvt  M31_5_ ( .D(net0115[2]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[2]));
nch_hvt  M31_4_ ( .D(net0115[3]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[3]));
nch_hvt  M31_3_ ( .D(net0115[4]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[4]));
nch_hvt  M31_2_ ( .D(net0115[5]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[5]));
nch_hvt  M31_1_ ( .D(net0115[6]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[6]));
nch_hvt  M31_0_ ( .D(net0115[7]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[7]));
nch_hvt  M19 ( .D(net0135), .B(GND_), .G(fsm_trim_ipp[0]),
     .S(net0131));
nch_hvt  M38_7_ ( .D(net0152[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_6_ ( .D(net0152[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_5_ ( .D(net0152[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_4_ ( .D(net0152[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_3_ ( .D(net0152[4]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_2_ ( .D(net0152[5]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_1_ ( .D(net0152[6]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_0_ ( .D(net0152[7]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_3_ ( .D(net0156[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_2_ ( .D(net0156[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_1_ ( .D(net0156[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_0_ ( .D(net0156[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_1_ ( .D(net0160[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_0_ ( .D(net0160[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M26 ( .D(net0131), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M33 ( .D(bl_pgm_glb), .B(GND_), .G(net0187), .S(gnd_));
nch_hvt  M30_3_ ( .D(net0172[0]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[0]));
nch_hvt  M30_2_ ( .D(net0172[1]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[1]));
nch_hvt  M30_1_ ( .D(net0172[2]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[2]));
nch_hvt  M30_0_ ( .D(net0172[3]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[3]));
nch_hvt  M34 ( .D(net089), .B(GND_), .G(pgm_trim0_en), .S(gnd_));
nch_hvt  M27_1_ ( .D(net0180[0]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[0]));
nch_hvt  M27_0_ ( .D(net0180[1]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[1]));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net0114), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net0114), .PLUS(net0141), .BULK(GND_));
inv_hvt I115 ( .A(net0116), .Y(net0187));
inv_hvt I58 ( .A(pgmen_b), .Y(pgmen));
inv_hvt I131 ( .A(fsm_pgm), .Y(pgmen_b));
inv_hvt I72 ( .A(fsm_pgmien_b_buf), .Y(fsm_pgmien_buf));
ml_ls_vdd2vdd25 I56 ( .in(pgmen), .sup(vddp_),
     .out_vddio_b(pgmen_b_25), .out_vddio(pgmen_25), .in_b(pgmen_b));
nch_25  M20 ( .D(net0173), .B(GND_), .G(pgm_inhi_bias),
     .S(bl_pgm_glb));
nch_25  M21 ( .D(pgm_inhi_bias), .B(GND_), .G(pgm_inhi_bias),
     .S(gnd_));
nch_25  M12_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[0]));
nch_25  M12_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[1]));
nch_25  M13_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[0]));
nch_25  M13_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[1]));
nch_25  M13_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[2]));
nch_25  M13_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[3]));
nch_25  M6 ( .D(net0164), .B(GND_), .G(net0164), .S(gnd_));
nch_25  M3 ( .D(dec_bias_p), .B(GND_), .G(bgr), .S(net0141));
nch_25  M10 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net089));
nch_25  M18_7_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[0]));
nch_25  M18_6_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[1]));
nch_25  M18_5_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[2]));
nch_25  M18_4_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[3]));
nch_25  M18_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[4]));
nch_25  M18_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[5]));
nch_25  M18_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[6]));
nch_25  M18_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[7]));
nch_25  M9 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net0135));
nch_25  M8 ( .D(net0164), .B(GND_), .G(pgmen_b_25), .S(gnd_));
pch_25  M11 ( .D(pgm_inhi_bias), .B(vddp_), .G(vdd_tieh), .S(net0259));
pch_25  M14_1_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M14_0_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M5 ( .D(net0164), .B(vddp_), .G(dec_bias_p), .S(net0199));
pch_25  M7_1_ ( .D(net0199), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M7_0_ ( .D(net0199), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M4 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p), .S(net0199));

endmodule
// Library - io, Cell - PDIDGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:24:26 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module PDIDGZ ( C, PAD );
output  C;

input  PAD;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_ymux_vblinhi_pgm_drv, View - schematic
// LAST TIME SAVED: Apr  8 10:44:07 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ymux_vblinhi_pgm_drv ( vblinhi_pgm_25, ysup_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25 );
inout  vblinhi_pgm_25, ysup_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd_), .B(GND_), .G(en_blinhi_pgm_b_ysup_25),
     .S(vblinhi_pgm_25));
pch_25  M5 ( .D(net10), .B(ysup_25), .G(en_blinhi_pgm_b_ysup_25),
     .S(ysup_25));
pch_25  M0 ( .D(net10), .B(vblinhi_pgm_25), .G(en_blinhi_pgm_b),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_wr_sup, View - schematic
// LAST TIME SAVED: Jan 24 10:11:13 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_wr_sup ( wr_sup_25, wrsup_2vdd, wrsup_2vdd_25 );
inout  wr_sup_25;

input  wrsup_2vdd, wrsup_2vdd_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I120 ( .A(net19), .Y(wrsup_vdd_in));
inv_hvt I131 ( .A(wrsup_2vdd), .Y(net19));
inv_25 I119 ( .IN(net20), .OUT(wrsup_vdd_in_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(wrsup_2vdd_25), .OUT(net20), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_2_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_1_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_0_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_ls25_1b, View - schematic
// LAST TIME SAVED: Jan 23 16:20:39 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25_1b ( out_25, in );
output  out_25;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I145 ( .A(in), .Y(net45));
inv_25 I153 ( .IN(out_b_25), .OUT(out_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I112 ( .in(in), .sup(vddp_), .out_vddio_b(out_b_25),
     .out_vddio(net025), .in_b(net45));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_ls25, View - schematic
// LAST TIME SAVED: May  1 10:33:06 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25 ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25,
     gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25, s_25,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wrsup_2vdd_25, fsm_gwlbdis, gnv, gred, gwl_misc, gwl_nvcm,
     gwl_red, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, s, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wrsup_2vdd_25;

input  fsm_gwlbdis, gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, testdec_en_b, testdec_even_b, testdec_odd_b,
     testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen, wrsup_2vdd;

output [5:0]  gnv_b_25;
output [3:0]  s_25;
output [1:0]  gred_25;
output [5:0]  gnv_25;
output [1:0]  gred_b_25;

input [5:0]  gnv;
input [3:0]  s;
input [1:0]  gred;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I_1_ ( .IN(gred_25[1]), .OUT(gred_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I_0_ ( .IN(gred_25[0]), .OUT(gred_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I143 ( .IN(net101), .OUT(fsm_gwlbdis_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_5_ ( .IN(gnv_25[5]), .OUT(gnv_b_25[5]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_4_ ( .IN(gnv_25[4]), .OUT(gnv_b_25[4]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_3_ ( .IN(gnv_25[3]), .OUT(gnv_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_2_ ( .IN(gnv_25[2]), .OUT(gnv_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_1_ ( .IN(gnv_25[1]), .OUT(gnv_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_0_ ( .IN(gnv_25[0]), .OUT(gnv_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_gwlwr_ctrl_ls25_1b I133 ( .in(testdec_en_b),
     .out_25(testdec_en_b_25));
ml_gwlwr_ctrl_ls25_1b I139 ( .in(gwlb_dis), .out_25(gwlb_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_frcen ( .in(wr_frcen),
     .out_25(wr_frcen_25));
ml_gwlwr_ctrl_ls25_1b I144 ( .in(gwlb_en), .out_25(gwlb_en_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vpp ( .in(gwphv_vppint),
     .out_25(gwphv_vppint_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwlb_vddp ( .in(gwlbsup_vddp),
     .out_25(gwlbsup_vddp_25));
ml_gwlwr_ctrl_ls25_1b ls25_gwlb_vpp ( .in(gwlbsup_vpxa),
     .out_25(gwlbsup_vpxa_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_vdd ( .in(wrsup_2vdd),
     .out_25(wrsup_2vdd_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_dis ( .in(wr_dis), .out_25(wr_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vddp ( .in(gwphv_vddp),
     .out_25(gwphv_vddp_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_frcen ( .in(wp_frcen),
     .out_25(wp_frcen_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_dis ( .in(wp_dis), .out_25(wp_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwl_red ( .in(gwl_red),
     .out_25(gwl_red_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_nvcm ( .in(gwl_nvcm),
     .out_25(gwl_nvcm_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_misc ( .in(gwl_misc),
     .out_25(gwl_misc_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_1_ ( .in(gred[1]),
     .out_25(gred_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_0_ ( .in(gred[0]),
     .out_25(gred_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_5_ ( .in(gnv[5]), .out_25(gnv_25[5]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_4_ ( .in(gnv[4]), .out_25(gnv_25[4]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_3_ ( .in(gnv[3]), .out_25(gnv_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_2_ ( .in(gnv[2]), .out_25(gnv_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_1_ ( .in(gnv[1]), .out_25(gnv_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_0_ ( .in(gnv[0]), .out_25(gnv_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_3_ ( .in(s[3]), .out_25(s_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_2_ ( .in(s[2]), .out_25(s_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_1_ ( .in(s[1]), .out_25(s_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_0_ ( .in(s[0]), .out_25(s_25[0]));
ml_gwlwr_ctrl_ls25_1b I134 ( .in(testdec_prec_b),
     .out_25(testdec_prec_b_25));
ml_gwlwr_ctrl_ls25_1b I136 ( .in(pgminhi_dmmy_b),
     .out_25(pgminhi_dmmy_b_25));
ml_gwlwr_ctrl_ls25_1b I140 ( .in(fsm_gwlbdis), .out_25(net101));
ml_gwlwr_ctrl_ls25_1b I137 ( .in(testdec_even_b),
     .out_25(testdec_even_b_25));
ml_gwlwr_ctrl_ls25_1b I138 ( .in(testdec_odd_b),
     .out_25(testdec_odd_b_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_npgate_gen, View - schematic
// LAST TIME SAVED: Sep 15 17:15:47 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa_npgate_gen ( dec_trim, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, vpxa, fsm_tm_testdec, saen, satrim,
     vddp_tieh );
output  saen_25, saen_b_vpxa;

inout  vpxa;

input  fsm_tm_testdec, saen, vddp_tieh;

output [4:1]  sa_ngate_25;
output [4:1]  sa_pgate_vpxa;
output [7:0]  dec_trim;

input [2:0]  satrim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net0122;

wire  [4:1]  trim_b;

wire  [4:1]  pgate_in;

wire  [7:0]  dec_trim_b;

wire  [0:3]  net48;

wire  [0:3]  net53;

wire  [4:1]  ngate_in_25_b;

wire  [2:0]  ydec_b;

wire  [2:0]  ydec;

wire  [4:1]  trim;



nor4_hvt I102 ( .D(fsm_tm_testdec), .C(dec_trim[7]), .A(dec_trim[5]),
     .B(dec_trim[6]), .Y(net47));
ml_hv_invx3 I135 ( .sel_hv(net048), .sel_25(net048),
     .vddp_tieh(vddp_tieh), .out_b_hv(saen_b_vpxa), .in_hv(vpxa));
ml_hv_invx3 I130_4_ ( .sel_hv(pgate_in[4]), .sel_25(pgate_in[4]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[4]), .in_hv(vpxa));
ml_hv_invx3 I130_3_ ( .sel_hv(pgate_in[3]), .sel_25(pgate_in[3]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[3]), .in_hv(vpxa));
ml_hv_invx3 I130_2_ ( .sel_hv(pgate_in[2]), .sel_25(pgate_in[2]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[2]), .in_hv(vpxa));
ml_hv_invx3 I130_1_ ( .sel_hv(pgate_in[1]), .sel_25(pgate_in[1]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[1]), .in_hv(vpxa));
inv_25 I149 ( .IN(net052), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I153_4_ ( .IN(ngate_in_25_b[4]), .OUT(sa_ngate_25[4]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_3_ ( .IN(ngate_in_25_b[3]), .OUT(sa_ngate_25[3]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_2_ ( .IN(ngate_in_25_b[2]), .OUT(sa_ngate_25[2]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_1_ ( .IN(ngate_in_25_b[1]), .OUT(sa_ngate_25[1]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_4_ ( .Y(dec_trim_b[4]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_3_ ( .Y(dec_trim_b[3]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_2_ ( .Y(dec_trim_b[2]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nand3_hvt I37_1_ ( .Y(dec_trim_b[1]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_0_ ( .Y(dec_trim_b[0]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nor2_hvt I75_4_ ( .Y(net48[0]), .B(dec_trim[4]), .A(sa_high_res));
nor2_hvt I75_3_ ( .Y(net48[1]), .B(dec_trim[3]), .A(trim[4]));
nor2_hvt I75_2_ ( .Y(net48[2]), .B(dec_trim[2]), .A(trim[3]));
nor2_hvt I75_1_ ( .Y(net48[3]), .B(dec_trim[1]), .A(trim[2]));
inv_hvt I145 ( .A(net076), .Y(net078));
inv_hvt I143 ( .A(net078), .Y(net080));
inv_hvt I146 ( .A(saen), .Y(net076));
inv_hvt I114 ( .A(net47), .Y(sa_high_res));
inv_hvt I38_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I38_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I38_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I38_4_ ( .A(dec_trim_b[4]), .Y(dec_trim[4]));
inv_hvt I38_3_ ( .A(dec_trim_b[3]), .Y(dec_trim[3]));
inv_hvt I38_2_ ( .A(dec_trim_b[2]), .Y(dec_trim[2]));
inv_hvt I38_1_ ( .A(dec_trim_b[1]), .Y(dec_trim[1]));
inv_hvt I38_0_ ( .A(dec_trim_b[0]), .Y(dec_trim[0]));
inv_hvt I40_2_ ( .A(ydec_b[2]), .Y(ydec[2]));
inv_hvt I40_1_ ( .A(ydec_b[1]), .Y(ydec[1]));
inv_hvt I40_0_ ( .A(ydec_b[0]), .Y(ydec[0]));
inv_hvt I76_4_ ( .A(net48[0]), .Y(trim[4]));
inv_hvt I76_3_ ( .A(net48[1]), .Y(trim[3]));
inv_hvt I76_2_ ( .A(net48[2]), .Y(trim[2]));
inv_hvt I76_1_ ( .A(net48[3]), .Y(trim[1]));
inv_hvt I39_2_ ( .A(satrim[2]), .Y(ydec_b[2]));
inv_hvt I39_1_ ( .A(satrim[1]), .Y(ydec_b[1]));
inv_hvt I39_0_ ( .A(satrim[0]), .Y(ydec_b[0]));
inv_hvt I78_4_ ( .A(trim[4]), .Y(trim_b[4]));
inv_hvt I78_3_ ( .A(trim[3]), .Y(trim_b[3]));
inv_hvt I78_2_ ( .A(trim[2]), .Y(trim_b[2]));
inv_hvt I78_1_ ( .A(trim[1]), .Y(trim_b[1]));
ml_ls_vdd2vdd25 I128_4_ ( .in(ngate_in_25_b[4]), .sup(vpxa),
     .out_vddio_b(pgate_in[4]), .out_vddio(net53[0]),
     .in_b(net0122[0]));
ml_ls_vdd2vdd25 I128_3_ ( .in(ngate_in_25_b[3]), .sup(vpxa),
     .out_vddio_b(pgate_in[3]), .out_vddio(net53[1]),
     .in_b(net0122[1]));
ml_ls_vdd2vdd25 I128_2_ ( .in(ngate_in_25_b[2]), .sup(vpxa),
     .out_vddio_b(pgate_in[2]), .out_vddio(net53[2]),
     .in_b(net0122[2]));
ml_ls_vdd2vdd25 I128_1_ ( .in(ngate_in_25_b[1]), .sup(vpxa),
     .out_vddio_b(pgate_in[1]), .out_vddio(net53[3]),
     .in_b(net0122[3]));
ml_ls_vdd2vdd25 I136 ( .in(net053), .sup(vpxa), .out_vddio_b(net047),
     .out_vddio(net048), .in_b(net052));
ml_ls_vdd2vdd25 I137 ( .in(net078), .sup(vddp_), .out_vddio_b(net052),
     .out_vddio(net053), .in_b(net080));
ml_ls_vdd2vdd25 I129_4_ ( .in(trim[4]), .sup(vddp_),
     .out_vddio_b(net0122[0]), .out_vddio(ngate_in_25_b[4]),
     .in_b(trim_b[4]));
ml_ls_vdd2vdd25 I129_3_ ( .in(trim[3]), .sup(vddp_),
     .out_vddio_b(net0122[1]), .out_vddio(ngate_in_25_b[3]),
     .in_b(trim_b[3]));
ml_ls_vdd2vdd25 I129_2_ ( .in(trim[2]), .sup(vddp_),
     .out_vddio_b(net0122[2]), .out_vddio(ngate_in_25_b[2]),
     .in_b(trim_b[2]));
ml_ls_vdd2vdd25 I129_1_ ( .in(trim[1]), .sup(vddp_),
     .out_vddio_b(net0122[3]), .out_vddio(ngate_in_25_b[1]),
     .in_b(trim_b[1]));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl, View - schematic
// LAST TIME SAVED: May  1 11:11:08 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25, gred_25,
     gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25,
     gwlb_en_25, pgminhi_dmmy_b_25, s_25, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv,
     vddp_tieh, vpp_int, vpxa, wr_sup_25, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

inout  bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv, vddp_tieh, vpp_int,
     vpxa, wr_sup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [5:0]  gnv_25;
output [5:0]  gnv_b_25;
output [1:0]  gred_25;
output [4:1]  sa_ngate_25;
output [3:0]  s_25;
output [1:0]  gred_b_25;
output [4:1]  sa_pgate_vpxa;

input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
input [0:0]  fsm_coladd;
input [3:0]  fsm_trim_ipp;
input [7:0]  fsm_rowadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  sa_trim;

wire  [3:0]  s;

wire  [1:0]  gred;

wire  [5:0]  gnv;

wire  [7:0]  dec_trim;



ml_hvmux_hotswitch_enhance Ihvmux_gwpsup_hv ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwphv_vppint_25), .sel_hv_a_25(gwphv_vddp_25),
     .out_hv(gwp_sup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_gwlwr_ctrl_logic Igwlwr_ctrl_logic ( .fsm_pgmdisc(fsm_pgmdisc),
     .gwlb_en(gwlb_en), .tm_testdec_wr(tm_testdec_wr),
     .tm_testdec(tm_testdec), .tm_dma(tm_dma),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_rd(fsm_rd), .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[0]), .wrsup_2vdd(wrsup_2vdd),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .testdec_prec_b(net172),
     .testdec_odd_b(testdec_odd_b), .testdec_even_b(testdec_even_b),
     .testdec_en_b(net175), .saen(saen), .sa_trim(sa_trim[2:0]),
     .s(s[3:0]), .pgminhi_dmmy_b(net179), .gwphv_vppint(gwphv_vppint),
     .gwphv_vddp(gwphv_vddp), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vddp(gwlbsup_vddp), .gwlb_dis(gwlb_dis),
     .gwl_misc(gwl_misc), .gred(gred[1:0]), .gnv(gnv[5:0]));
ml_hvmux_hotswitch Ihvmux_gwlbsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwlbsup_vpxa_25), .sel_hv_a_25(gwlbsup_vddp_25),
     .out_hv(gwl_b_sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_gwlwr_bldrv Igwlwr_bldrv ( .fsm_din(fsm_din), .tm_dma(tm_dma),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .bl_frc_gnd(gnd_), .bgr(bgr),
     .bl_pgm_glb(bl_pgm_glb));
ml_gwlwr_ctrl_wr_sup Igwlwr_ctrl_wr_sup ( .wrsup_2vdd(wrsup_2vdd),
     .wrsup_2vdd_25(wrsup_2vdd_25), .wr_sup_25(wr_sup_25));
ml_gwlwr_ctrl_ls25 Igwlwr_ctrl_ls25 ( .gwlb_en_25(gwlb_en_25),
     .gwlb_en(gwlb_en), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwlb_dis(gwlb_dis), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vpxa_25(gwlbsup_vpxa_25), .wrsup_2vdd_25(wrsup_2vdd_25),
     .wrsup_2vdd(wrsup_2vdd), .testdec_odd_b(testdec_odd_b),
     .testdec_even_b(testdec_even_b),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .testdec_prec_b(net172),
     .testdec_en_b(net175), .pgminhi_dmmy_b(net179),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwphv_vddp(gwphv_vddp),
     .gwlbsup_vddp(gwlbsup_vddp), .gwphv_vppint(gwphv_vppint),
     .gwlbsup_vddp_25(gwlbsup_vddp_25),
     .gwphv_vppint_25(gwphv_vppint_25), .gwphv_vddp_25(gwphv_vddp_25),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .s(s[3:0]), .gwl_red(fsm_nv_rrow),
     .gwl_nvcm(fsm_nv_bstream), .gwl_misc(gwl_misc), .gred(gred[1:0]),
     .gnv(gnv[5:0]), .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]));
vddp_tiehigh Ivddp_tiehigh_15_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_14_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_13_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_12_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_11_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_10_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_9_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_8_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_0_ ( .vddp_tieh(vddp_tieh));
ml_core_sa_npgate_gen Icore_sa_npgate_gen (
     .fsm_tm_testdec(tm_testdec), .satrim(sa_trim[2:0]),
     .vddp_tieh(vddp_tieh), .saen(saen), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .dec_trim(dec_trim[7:0]),
     .vpxa(vpxa));

endmodule
// Library - NVCM, Cell - ml_gwlwr_top_1f, View - schematic
// LAST TIME SAVED: Jan 20 17:29:58 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_gwlwr_top_1f ( fsm_gwlbdis_b_25, gwl_b_25, gwl_b_sup_25,
     gwp_hv, pgminhi_dmmy_b_25, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wr, bgr, bl_pgm_glb, vpp_int, vpxa, fsm_coladd,
     fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_b_sup_25, pgminhi_dmmy_b_25, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25;

inout  bgr, bl_pgm_glb, vpp_int, vpxa;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [26:0]  gwp_hv;
output [4:1]  sa_ngate_25;
output [4:1]  sa_pgate_vpxa;
output [26:0]  gwl_b_25;
output [107:0]  wr;

input [2:0]  fsm_trim_rrefrd;
input [7:0]  fsm_rowadd;
input [0:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_trim_ipp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  gnv_25;

wire  [5:0]  gnv_b_25;

wire  [1:0]  gred_25;

wire  [1:0]  gred_b_25;

wire  [3:0]  s_25;



ml_gwlwr_1f Igwlwr_1f ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .gwlb_en_25(gwlb_en_25), .gwlb_dis_25(gwlb_dis_25),
     .wr_sup_25(wr_sup_25), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .vddp_tieh(vddp_tieh), .s_25(s_25[3:0]),
     .gwl_red_25(gwl_red_25), .gwl_nvcm_25(gwl_nvcm_25),
     .gwl_misc_25(gwl_misc_25), .gred_b_25(gred_b_25[1:0]),
     .gred_25(gred_25[1:0]), .gnv_b_25(gnv_b_25[5:0]),
     .gnv_25(gnv_25[5:0]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25));
ml_gwlwr_ctrl Igwlwr_ctrl ( .fsm_pgmdisc(fsm_pgmdisc),
     .gwlb_en_25(gwlb_en_25), .fsm_din(fsm_din),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_allwl_l(fsm_tm_allwl_l), .fsm_tm_allwl_h(fsm_tm_allwl_h),
     .fsm_tm_allbl_l(fsm_tm_allbl_l), .fsm_tm_allbl_h(fsm_tm_allbl_h),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .s_25(s_25[3:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwl_red_25(gwl_red_25), .gwl_nvcm_25(gwl_nvcm_25),
     .gwl_misc_25(gwl_misc_25), .gred_b_25(gred_b_25[1:0]),
     .gred_25(gred_25[1:0]), .gnv_b_25(gnv_b_25[5:0]),
     .gnv_25(gnv_25[5:0]), .wr_sup_25(wr_sup_25), .vpxa(vpxa),
     .vpp_int(vpp_int), .vddp_tieh(vddp_tieh), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr));

endmodule
// Library - NVCM, Cell - ml_core_sa_spare, View - schematic
// LAST TIME SAVED: Sep 22 17:28:46 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa_spare (  );supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:9]  net501;



rppolywo_m  R7 ( .MINUS(net033), .PLUS(net036), .BULK(gnd_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(net033), .BULK(gnd_));
rppolywo_m  R3 ( .MINUS(net042), .PLUS(net039), .BULK(gnd_));
rppolywo_m  R4 ( .MINUS(gnd_), .PLUS(net042), .BULK(gnd_));
rppolywo_m  R5 ( .MINUS(net039), .PLUS(net045), .BULK(gnd_));
rppolywo_m  R6 ( .MINUS(net045), .PLUS(net027), .BULK(gnd_));
rppolywo_m  R9 ( .MINUS(net036), .PLUS(net030), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(net030), .PLUS(net027), .BULK(gnd_));
vdd_tielow I144_9_ ( .gnd_tiel(net501[0]));
vdd_tielow I144_8_ ( .gnd_tiel(net501[1]));
vdd_tielow I144_7_ ( .gnd_tiel(net501[2]));
vdd_tielow I144_6_ ( .gnd_tiel(net501[3]));
vdd_tielow I144_5_ ( .gnd_tiel(net501[4]));
vdd_tielow I144_4_ ( .gnd_tiel(net501[5]));
vdd_tielow I144_3_ ( .gnd_tiel(net501[6]));
vdd_tielow I144_2_ ( .gnd_tiel(net501[7]));
vdd_tielow I144_1_ ( .gnd_tiel(net501[8]));
vdd_tielow I144_0_ ( .gnd_tiel(net501[9]));

endmodule
// Library - NVCM, Cell - ml_testdec_rows, View - schematic
// LAST TIME SAVED: Feb 26 14:35:11 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_testdec_rows ( dec_bias, dec_det_25, vddp_tieh, wp, wr );
inout  dec_bias, dec_det_25;

input  vddp_tieh, wp, wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(dec_det_25), .B(GND_), .G(wr), .S(gnd_));
nch_25  M12 ( .D(net20), .B(gnd_), .G(vddp_tieh), .S(wp));
nch_25  M2 ( .D(dec_det_25), .B(GND_), .G(net20), .S(gnd_));
nch_25  M0 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(net20));
nch_25  M1 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(wr));

endmodule
// Library - NVCM, Cell - ml_testdec_rowsx108_1f, View - schematic
// LAST TIME SAVED: Jan 20 11:17:22 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_testdec_rowsx108_1f ( dec_det_even_25, dec_det_odd_25,
     dec_bias_25, dec_det_25, testdec_even_b_25, testdec_odd_b_25, wp,
     wr );
output  dec_det_even_25, dec_det_odd_25;

inout  dec_bias_25, dec_det_25;

input  testdec_even_b_25, testdec_odd_b_25;

input [107:0]  wr;
input [107:0]  wp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I25 ( .vddp_tieh(vddp_tiel));
nor2_25 I24 ( .A(testdec_odd_b_25), .Y(dec_det_odd_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
nor2_25 I59 ( .A(testdec_even_b_25), .Y(dec_det_even_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
ml_testdec_rows Itestdec_rows_107_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[107]), .wp(wp[107]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_106_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[106]), .wp(wp[106]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_105_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[105]), .wp(wp[105]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_104_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[104]), .wp(wp[104]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_103_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[103]), .wp(wp[103]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_102_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[102]), .wp(wp[102]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_101_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[101]), .wp(wp[101]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_100_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[100]), .wp(wp[100]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_99_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[99]), .wp(wp[99]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_98_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[98]), .wp(wp[98]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_97_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[97]), .wp(wp[97]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_96_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[96]), .wp(wp[96]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_95_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[95]), .wp(wp[95]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_94_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[94]), .wp(wp[94]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_93_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[93]), .wp(wp[93]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_92_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[92]), .wp(wp[92]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_91_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[91]), .wp(wp[91]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_90_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[90]), .wp(wp[90]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_89_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[89]), .wp(wp[89]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_88_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[88]), .wp(wp[88]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_87_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[87]), .wp(wp[87]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_86_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[86]), .wp(wp[86]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_85_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[85]), .wp(wp[85]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_84_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[84]), .wp(wp[84]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_83_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[83]), .wp(wp[83]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_82_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[82]), .wp(wp[82]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_81_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[81]), .wp(wp[81]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_80_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[80]), .wp(wp[80]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_79_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[79]), .wp(wp[79]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_78_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[78]), .wp(wp[78]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_77_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[77]), .wp(wp[77]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_76_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[76]), .wp(wp[76]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_75_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[75]), .wp(wp[75]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_74_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[74]), .wp(wp[74]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_73_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[73]), .wp(wp[73]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_72_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[72]), .wp(wp[72]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_71_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[71]), .wp(wp[71]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_70_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[70]), .wp(wp[70]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_69_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[69]), .wp(wp[69]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_68_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[68]), .wp(wp[68]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_67_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[67]), .wp(wp[67]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_66_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[66]), .wp(wp[66]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_65_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[65]), .wp(wp[65]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_64_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[64]), .wp(wp[64]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_63_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[63]), .wp(wp[63]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_62_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[62]), .wp(wp[62]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_61_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[61]), .wp(wp[61]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_60_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[60]), .wp(wp[60]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_59_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[59]), .wp(wp[59]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_58_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[58]), .wp(wp[58]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_57_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[57]), .wp(wp[57]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_56_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[56]), .wp(wp[56]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_55_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[55]), .wp(wp[55]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_54_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[54]), .wp(wp[54]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_53_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[53]), .wp(wp[53]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_52_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[52]), .wp(wp[52]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_51_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[51]), .wp(wp[51]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_50_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[50]), .wp(wp[50]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_49_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[49]), .wp(wp[49]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_48_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[48]), .wp(wp[48]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_47_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[47]), .wp(wp[47]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_46_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[46]), .wp(wp[46]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_45_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[45]), .wp(wp[45]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_44_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[44]), .wp(wp[44]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_43_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[43]), .wp(wp[43]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_42_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[42]), .wp(wp[42]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_41_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[41]), .wp(wp[41]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_40_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[40]), .wp(wp[40]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_39_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[39]), .wp(wp[39]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_38_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[38]), .wp(wp[38]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_37_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[37]), .wp(wp[37]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_36_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[36]), .wp(wp[36]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_35_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[35]), .wp(wp[35]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_34_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[34]), .wp(wp[34]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_33_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[33]), .wp(wp[33]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_32_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[32]), .wp(wp[32]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_31_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[31]), .wp(wp[31]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_30_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[30]), .wp(wp[30]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_29_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[29]), .wp(wp[29]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_28_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[28]), .wp(wp[28]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_27_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[27]), .wp(wp[27]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_26_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[26]), .wp(wp[26]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_25_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[25]), .wp(wp[25]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_24_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[24]), .wp(wp[24]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_23_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[23]), .wp(wp[23]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_22_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[22]), .wp(wp[22]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_21_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[21]), .wp(wp[21]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_20_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[20]), .wp(wp[20]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_19_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[19]), .wp(wp[19]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_18_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[18]), .wp(wp[18]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_17_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[17]), .wp(wp[17]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_16_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[16]), .wp(wp[16]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_15_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[15]), .wp(wp[15]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_14_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[14]), .wp(wp[14]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_13_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[13]), .wp(wp[13]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_12_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[12]), .wp(wp[12]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_11_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[11]), .wp(wp[11]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_10_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[10]), .wp(wp[10]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_9_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[9]), .wp(wp[9]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_8_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[8]), .wp(wp[8]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_7_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[7]), .wp(wp[7]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_6_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[6]), .wp(wp[6]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_5_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[5]), .wp(wp[5]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_4_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[4]), .wp(wp[4]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_3_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[3]), .wp(wp[3]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_2_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[2]), .wp(wp[2]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_1_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[1]), .wp(wp[1]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_0_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[0]), .wp(wp[0]),
     .dec_bias(dec_bias_25));

endmodule
// Library - io, Cell - PDU08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 17:45:09 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module PDU08DGZ ( C, PAD, I, OEN );
output  C;

inout  PAD;

input  I, OEN;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_rock_gwlgnd_nor2, View - schematic
// LAST TIME SAVED: Jan 23 10:17:03 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_rock_gwlgnd_nor2 ( gwl_gnd_25, gwl_b_sup_25, gwl_b_25,
     gwl_b_gnden_25 );
output  gwl_gnd_25;

inout  gwl_b_sup_25;

input  gwl_b_25, gwl_b_gnden_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(net14), .B(GND_), .G(gwl_b_gnden_25), .S(GND_));
nch_25  M0 ( .D(gwl_gnd_25), .B(GND_), .G(gwl_b_25), .S(net14));
pch_25  M2 ( .D(gwl_gnd_25), .B(gwl_b_sup_25), .G(gwl_b_25),
     .S(gwl_b_sup_25));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp, View - schematic
// LAST TIME SAVED: Jan 21 10:22:42 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp ( wp, ngate_25, gwl_b_25, gwl_gnd_25, gwp_hv,
     s_b_25, s_b_hv );
output  wp;

inout  ngate_25;

input  gwl_b_25, gwl_gnd_25, gwp_hv, s_b_25, s_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M6 ( .D(wp), .B(gwp_hv), .G(s_b_hv), .S(gwp_hv));
nch_25  M11 ( .D(net18), .B(GND_), .G(s_b_25), .S(gwl_gnd_25));
nch_25  M12 ( .D(wp), .B(GND_), .G(ngate_25), .S(net18));
nch_25  M10 ( .D(net18), .B(GND_), .G(gwl_b_25), .S(gwl_gnd_25));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp_x4, View - schematic
// LAST TIME SAVED: Jan 23 10:17:05 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x4 ( wp, gwl_b_sup_25, ngate_25, gwl_b_25,
     gwl_b_gnden_25, gwp_hv, s_b_25, s_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_25, gwl_b_gnden_25, gwp_hv;

output [3:0]  wp;

input [3:0]  s_b_25;
input [3:0]  s_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwl_b_25(gwl_b_25), .gwl_gnd_25(gwl_gnd_25));
ml_rock_lwldrv_wp Iml_lwldrv_1 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[1]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[1]), .wp(wp[1]));
ml_rock_lwldrv_wp Iml_lwldrv_2 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[2]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[2]), .wp(wp[2]));
ml_rock_lwldrv_wp Iml_lwldrv_3 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[3]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3]), .wp(wp[3]));
ml_rock_lwldrv_wp Iml_lwldrv_0 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[0]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[0]), .wp(wp[0]));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp_x108_1f, View - schematic
// LAST TIME SAVED: Jan 20 11:13:16 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x108_1f ( wp, gwl_b_sup_25, ngate_25, s_b_25,
     s_b_hv, gwl_b_25, gwl_b_gnden_25, gwp_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_gnden_25;

output [107:0]  wp;

inout [3:0]  s_b_25;
inout [3:0]  s_b_hv;

input [26:0]  gwl_b_25;
input [26:0]  gwp_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_26_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[26]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[107:104]), .gwl_b_25(gwl_b_25[26]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_25_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[25]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[103:100]), .gwl_b_25(gwl_b_25[25]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_24_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[24]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[99:96]), .gwl_b_25(gwl_b_25[24]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_23_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[23]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[95:92]), .gwl_b_25(gwl_b_25[23]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_22_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[22]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[91:88]), .gwl_b_25(gwl_b_25[22]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_21_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[21]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[87:84]), .gwl_b_25(gwl_b_25[21]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_20_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[20]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[83:80]), .gwl_b_25(gwl_b_25[20]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_19_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[19]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[79:76]), .gwl_b_25(gwl_b_25[19]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_18_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[18]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[75:72]), .gwl_b_25(gwl_b_25[18]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_17_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[17]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[71:68]), .gwl_b_25(gwl_b_25[17]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_16_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[16]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[67:64]), .gwl_b_25(gwl_b_25[16]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_15_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[15]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[63:60]), .gwl_b_25(gwl_b_25[15]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_14_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[14]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[59:56]), .gwl_b_25(gwl_b_25[14]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_13_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[13]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[55:52]), .gwl_b_25(gwl_b_25[13]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_12_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[12]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[51:48]), .gwl_b_25(gwl_b_25[12]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_11_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[11]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[47:44]), .gwl_b_25(gwl_b_25[11]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_10_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[10]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[43:40]), .gwl_b_25(gwl_b_25[10]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_9_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[9]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[39:36]), .gwl_b_25(gwl_b_25[9]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_8_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[8]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[35:32]), .gwl_b_25(gwl_b_25[8]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_7_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[7]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[31:28]), .gwl_b_25(gwl_b_25[7]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_6_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[6]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[27:24]), .gwl_b_25(gwl_b_25[6]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_5_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[5]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[23:20]), .gwl_b_25(gwl_b_25[5]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_4_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[4]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[19:16]), .gwl_b_25(gwl_b_25[4]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_3_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[3]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[15:12]), .gwl_b_25(gwl_b_25[3]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_2_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[2]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[11:8]), .gwl_b_25(gwl_b_25[2]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_1_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[1]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[7:4]), .gwl_b_25(gwl_b_25[1]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_0_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[0]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[3:0]), .gwl_b_25(gwl_b_25[0]), .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - ROCK, Cell - nvcm_cell_1, View - schematic
// LAST TIME SAVED: May 13 16:00:35 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module nvcm_cell_1 ( bl, wp, wr );
inout  bl;

input  wp, wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nchx  NR ( .D(net1), .G(wr), .S(bl));
nchx  NP ( .D(net5), .G(wp), .S(net1));

endmodule
// Library - NVCM, Cell - nvcm_cell_2x1, View - schematic
// LAST TIME SAVED: Dec 10 15:56:30 2007
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module nvcm_cell_2x1 ( bl, wp, wr );

input  wp, wr;

inout [1:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
nvcm_cell_1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));

endmodule
// Library - NVCM, Cell - nvcm_cell_2x8, View - schematic
// LAST TIME SAVED: Feb 26 14:36:29 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module nvcm_cell_2x8 ( bl, wp, wr );


inout [1:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x1 m7 ( .bl(bl[1:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_2x1 m6 ( .bl(bl[1:0]), .wr(wr[6]), .wp(wp[6]));
nvcm_cell_2x1 m5 ( .bl(bl[1:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_2x1 m4 ( .bl(bl[1:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_2x1 m3 ( .bl(bl[1:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_2x1 m2 ( .bl(bl[1:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_2x1 m1 ( .bl(bl[1:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_2x1 m0 ( .bl(bl[1:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM, Cell - nvcm_cell_1x8, View - schematic
// LAST TIME SAVED: Jul  5 11:06:02 2007
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module nvcm_cell_1x8 ( bl, wp, wr );

input  wp, wr;

inout [7:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
nvcm_cell_1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));
nvcm_cell_1 m2 ( .wp(wp), .wr(wr), .bl(bl[2]));
nvcm_cell_1 m3 ( .wp(wp), .wr(wr), .bl(bl[3]));
nvcm_cell_1 m4 ( .wp(wp), .wr(wr), .bl(bl[4]));
nvcm_cell_1 m5 ( .wp(wp), .wr(wr), .bl(bl[5]));
nvcm_cell_1 m6 ( .wp(wp), .wr(wr), .bl(bl[6]));
nvcm_cell_1 m7 ( .wp(wp), .wr(wr), .bl(bl[7]));

endmodule
// Library - NVCM, Cell - nvcm_cell_8x8, View - schematic
// LAST TIME SAVED: Dec 10 15:35:50 2007
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module nvcm_cell_8x8 ( bl, wp, wr );


inout [7:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1x8 m0 ( .bl(bl[7:0]), .wr(wr[0]), .wp(wp[0]));
nvcm_cell_1x8 m1 ( .bl(bl[7:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 m2 ( .bl(bl[7:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_1x8 m3 ( .bl(bl[7:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_1x8 m7 ( .bl(bl[7:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_1x8 m4 ( .bl(bl[7:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_1x8 m5 ( .bl(bl[7:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_1x8 m6 ( .bl(bl[7:0]), .wr(wr[6]), .wp(wp[6]));

endmodule
// Library - NVCM, Cell - nvcm_cell_16x8, View - schematic
// LAST TIME SAVED: Dec 10 15:41:25 2007
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module nvcm_cell_16x8 ( bl, wp, wr );


inout [15:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_8x8 m0 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[7:0]));
nvcm_cell_8x8 m1 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[15:8]));

endmodule
// Library - io, Cell - botbank_1k_july16, View - schematic
// LAST TIME SAVED: Jul 16 12:54:14 2009
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module botbank_1k_july16 ( cdone_int, ctst_b_int, in, done, pad,
     cdone_out, ctst_b, oen, out, ren );
output  cdone_int, ctst_b_int;

inout  done;

input  cdone_out, ctst_b;

output [23:0]  in;

inout [23:0]  pad;

input [23:0]  oen;
input [23:0]  out;
input [23:0]  ren;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



PVDD1DGZ I76_1_ ( .VDD(vdd_));
PVDD1DGZ I76_0_ ( .VDD(vdd_));
PDIDGZ I41 ( .PAD(ctst_b), .C(ctst_b_int));
PDU08DGZ I39 ( .PAD(done), .C(cdone_int), .OEN(cdone_out), .I(gnd_));
PDUW08DGZ I72_21_ ( .PAD(pad[21]), .C(in[21]), .OEN(oen[21]),
     .I(out[21]), .REN(ren[21]));
PDUW08DGZ I72_20_ ( .PAD(pad[20]), .C(in[20]), .OEN(oen[20]),
     .I(out[20]), .REN(ren[20]));
PDUW08DGZ I77_19_ ( .PAD(pad[19]), .C(in[19]), .OEN(oen[19]),
     .I(out[19]), .REN(ren[19]));
PDUW08DGZ I77_18_ ( .PAD(pad[18]), .C(in[18]), .OEN(oen[18]),
     .I(out[18]), .REN(ren[18]));
PDUW08DGZ I77_17_ ( .PAD(pad[17]), .C(in[17]), .OEN(oen[17]),
     .I(out[17]), .REN(ren[17]));
PDUW08DGZ I77_16_ ( .PAD(pad[16]), .C(in[16]), .OEN(oen[16]),
     .I(out[16]), .REN(ren[16]));
PDUW08DGZ I77_15_ ( .PAD(pad[15]), .C(in[15]), .OEN(oen[15]),
     .I(out[15]), .REN(ren[15]));
PDUW08DGZ I40_9_ ( .PAD(pad[9]), .C(in[9]), .OEN(oen[9]), .I(out[9]),
     .REN(ren[9]));
PDUW08DGZ I40_8_ ( .PAD(pad[8]), .C(in[8]), .OEN(oen[8]), .I(out[8]),
     .REN(ren[8]));
PDUW08DGZ I67_7_ ( .PAD(pad[7]), .C(in[7]), .OEN(oen[7]), .I(out[7]),
     .REN(ren[7]));
PDUW08DGZ I67_6_ ( .PAD(pad[6]), .C(in[6]), .OEN(oen[6]), .I(out[6]),
     .REN(ren[6]));
PDUW08DGZ I67_5_ ( .PAD(pad[5]), .C(in[5]), .OEN(oen[5]), .I(out[5]),
     .REN(ren[5]));
PDUW08DGZ I67_4_ ( .PAD(pad[4]), .C(in[4]), .OEN(oen[4]), .I(out[4]),
     .REN(ren[4]));
PDUW08DGZ I67_3_ ( .PAD(pad[3]), .C(in[3]), .OEN(oen[3]), .I(out[3]),
     .REN(ren[3]));
PDUW08DGZ I67_2_ ( .PAD(pad[2]), .C(in[2]), .OEN(oen[2]), .I(out[2]),
     .REN(ren[2]));
PDUW08DGZ I67_1_ ( .PAD(pad[1]), .C(in[1]), .OEN(oen[1]), .I(out[1]),
     .REN(ren[1]));
PDUW08DGZ I67_0_ ( .PAD(pad[0]), .C(in[0]), .OEN(oen[0]), .I(out[0]),
     .REN(ren[0]));
PDUW08DGZ I43_23_ ( .PAD(pad[23]), .C(in[23]), .OEN(oen[23]),
     .I(out[23]), .REN(ren[23]));
PDUW08DGZ I43_22_ ( .PAD(pad[22]), .C(in[22]), .OEN(oen[22]),
     .I(out[22]), .REN(ren[22]));
PDUW08DGZ I75_11_ ( .PAD(pad[11]), .C(in[11]), .OEN(oen[11]),
     .I(out[11]), .REN(ren[11]));
PDUW08DGZ I75_10_ ( .PAD(pad[10]), .C(in[10]), .OEN(oen[10]),
     .I(out[10]), .REN(ren[10]));
PDUW08DGZ I66_13_ ( .PAD(pad[13]), .C(in[13]), .OEN(oen[13]),
     .I(out[13]), .REN(ren[13]));
PDUW08DGZ I66_12_ ( .PAD(pad[12]), .C(in[12]), .OEN(oen[12]),
     .I(out[12]), .REN(ren[12]));
PDUW08DGZ I68_14_ ( .PAD(pad[14]), .C(in[14]), .OEN(oen[14]),
     .I(out[14]), .REN(ren[14]));
PVDD2DGZ I56 ( .VDDPST(vddio_spi));
PVDD2DGZ I74_1_ ( .VDDPST(vddio_bottombank));
PVDD2DGZ I74_0_ ( .VDDPST(vddio_bottombank));
PVDD2DGZ I69_1_ ( .VDDPST(vddio_bottombank));
PVDD2DGZ I69_0_ ( .VDDPST(vddio_bottombank));
PVDD2POC I57 ( .VDDPST(vddio_spi));
PVDD2POC I71 ( .VDDPST(vddio_bottombank));
PVSS3DGZ I62_1_ ( .VSS(gnd_));
PVSS3DGZ I62_0_ ( .VSS(gnd_));
PVSS3DGZ I73_1_ ( .VSS(gnd_));
PVSS3DGZ I73_0_ ( .VSS(gnd_));
PVSS3DGZ I64_2_ ( .VSS(gnd_));
PVSS3DGZ I64_1_ ( .VSS(gnd_));
PVSS3DGZ I64_0_ ( .VSS(gnd_));

endmodule
// Library - NVCM, Cell - nvcm_cell_336x8, View - schematic
// LAST TIME SAVED: Feb 26 14:32:20 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module nvcm_cell_336x8 ( bl, bl_dummyl, bl_dummyr, bl_test, wp, wr );


inout [1:0]  bl_test;
inout [327:0]  bl;
inout [1:0]  bl_dummyl;
inout [5:0]  bl_dummyr;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x8 Invcm_cell_2x8 ( .wp(wp[7:0]), .wr(wr[7:0]),
     .bl(bl_dummyl[1:0]));
nvcm_cell_16x8 Invcm_cell_16x8_19_ ( .wp(wp[7:0]), .bl(bl[319:304]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_18_ ( .wp(wp[7:0]), .bl(bl[303:288]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_17_ ( .wp(wp[7:0]), .bl(bl[287:272]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_16_ ( .wp(wp[7:0]), .bl(bl[271:256]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_15_ ( .wp(wp[7:0]), .bl(bl[255:240]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_14_ ( .wp(wp[7:0]), .bl(bl[239:224]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_13_ ( .wp(wp[7:0]), .bl(bl[223:208]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_12_ ( .wp(wp[7:0]), .bl(bl[207:192]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_11_ ( .wp(wp[7:0]), .bl(bl[191:176]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_10_ ( .wp(wp[7:0]), .bl(bl[175:160]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_9_ ( .wp(wp[7:0]), .bl(bl[159:144]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_8_ ( .wp(wp[7:0]), .bl(bl[143:128]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_7_ ( .wp(wp[7:0]), .bl(bl[127:112]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_6_ ( .wp(wp[7:0]), .bl(bl[111:96]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_5_ ( .wp(wp[7:0]), .bl(bl[95:80]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_4_ ( .wp(wp[7:0]), .bl(bl[79:64]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_3_ ( .wp(wp[7:0]), .bl(bl[63:48]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_2_ ( .wp(wp[7:0]), .bl(bl[47:32]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_1_ ( .wp(wp[7:0]), .bl(bl[31:16]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_0_ ( .wp(wp[7:0]), .bl(bl[15:0]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_20_ ( .wp(wp[7:0]), .bl({bl_dummyr[5:0],
     bl_test[1:0], bl[327:320]}), .wr(wr[7:0]));

endmodule
// Library - NVCM, Cell - nvcm_cell_338x112_1f, View - schematic
// LAST TIME SAVED: Jan 20 11:01:43 2009
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module nvcm_cell_338x112_1f ( bl, bl_dummyl, bl_dummyr, bl_test, wp,
     wp_dummyb, wp_dummyt, wr, wr_dummyb, wr_dummyt );


inout [327:0]  bl;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;
inout [1:0]  bl_dummyr;

input [1:0]  wp_dummyt;
input [1:0]  wr_dummyb;
input [1:0]  wp_dummyb;
input [107:0]  wp;
input [1:0]  wr_dummyt;
input [107:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_336x8 Invcm_cell_336x8_11_ ( .wr(wr[101:94]),
     .wp(wp[101:94]), .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_10_ ( .wr(wr[93:86]), .wp(wp[93:86]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_9_ ( .wr(wr[85:78]), .wp(wp[85:78]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_8_ ( .wr(wr[77:70]), .wp(wp[77:70]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_7_ ( .wr(wr[69:62]), .wp(wp[69:62]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_6_ ( .wr(wr[61:54]), .wp(wp[61:54]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_5_ ( .wr(wr[53:46]), .wp(wp[53:46]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_4_ ( .wr(wr[45:38]), .wp(wp[45:38]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_3_ ( .wr(wr[37:30]), .wp(wp[37:30]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_2_ ( .wr(wr[29:22]), .wp(wp[29:22]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_1_ ( .wr(wr[21:14]), .wp(wp[21:14]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_0_ ( .wr(wr[13:6]), .wp(wp[13:6]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_t ( .wr({wr[5:0], wr_dummyt[1:0]}),
     .wp({wp[5:0], wp_dummyt[1:0]}), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_b ( .wr({wr_dummyb[1:0],
     wr[107:102]}), .wp({wp_dummyb[1:0], wp[107:102]}),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));

endmodule
// Library - sbtlibn65lp, Cell - oai221x2_hvt, View - schematic
// LAST TIME SAVED: May  4 14:29:05 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module oai221x2_hvt ( Y, A0, A1, B0, B1, C0 );
output  Y;

input  A0, A1, B0, B1, C0;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(net040), .B(GND_), .G(A0), .S(net024));
nch_hvt  M11 ( .D(Y), .B(GND_), .G(C0), .S(net040));
nch_hvt  M8 ( .D(net040), .B(GND_), .G(A1), .S(net024));
nch_hvt  M10 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
pch_hvt  M7 ( .D(Y), .B(VDD_), .G(C0), .S(vdd_));
pch_hvt  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M4 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
pch_hvt  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_ls_vdd25_nor2, View - schematic
// LAST TIME SAVED: Jan 12 15:33:21 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_ls_vdd25_nor2 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_25 I79 ( .A(in), .Y(out_vddio_b), .Gb(gnd_), .G(gnd_), .Pb(sup),
     .P(sup), .B(out_vddio));
nor2_25 I151 ( .A(out_vddio_b), .Y(out_vddio), .Gb(gnd_), .G(gnd_),
     .Pb(sup), .P(sup), .B(in_b));

endmodule
// Library - NVCM, Cell - ml_core_ctrl_logic, View - schematic
// LAST TIME SAVED: May 12 10:24:23 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_ctrl_logic ( dec_trim, en_blinhi_pgm_b,
     en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25, yp1_sel,
     yp2_sel, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, yp21_b_low_b, yp_test, fsm_blkadd,
     fsm_coladd, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, tm_tcol, ysup_25 );
output  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp21_b_low_b;

input  fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h,
     fsm_tm_allwl_l, fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, tm_tcol, ysup_25;

output [7:0]  yp3_sel;
output [3:0]  sb25_high_25;
output [3:0]  sbhv_high_25;
output [3:0]  sb25_gnd_25;
output [7:0]  yp2_sel;
output [1:0]  yp_test;
output [7:5]  dec_trim;
output [5:0]  yp1_sel;
output [3:0]  sbhv_gnd_25;

input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefpgm;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net319;

wire  [7:0]  yp2_sel_b;

wire  [7:0]  yp3_sel_b;

wire  [7:5]  dec_trim_b;

wire  [2:0]  tdec_b;

wire  [2:0]  tdec;

wire  [3:0]  sb25low_b;

wire  [1:0]  yp_test_b;

wire  [0:3]  net339;

wire  [0:3]  net317;

wire  [1:0]  xadd;

wire  [3:0]  sbhvlow_b;

wire  [1:0]  xadd_b;

wire  [5:0]  yp1_sel_b;

wire  [8:0]  yadd;

wire  [8:0]  yadd_b;

wire  [0:3]  net387;

wire  [0:3]  net523;

wire  [0:3]  net407;

wire  [0:3]  net299;

wire  [0:3]  net522;

wire  [0:3]  net323;

wire  [0:3]  net393;

wire  [0:3]  net409;

wire  [0:3]  net304;

wire  [0:3]  net552;

wire  [0:3]  net546;

wire  [0:3]  net321;

wire  [0:2]  net629;

wire  [0:3]  net411;

wire  [0:3]  net391;

wire  [0:3]  net549;

wire  [0:3]  net544;



oai21x2 I36 ( .A1(fsm_pgmvfy), .A0(fsm_rd), .B0(net425),
     .Y(all_blk_sel_b));
oai221x2_hvt I86_3_ ( .C0(yadd_b[8]), .A1(net565), .Y(yp1_sel_b[3]),
     .A0(yadd[7]), .B0(vddp_rd_overw), .B1(yadd[6]));
oai221x2_hvt I86_2_ ( .C0(yadd_b[8]), .A1(net565), .Y(yp1_sel_b[2]),
     .A0(yadd[7]), .B0(vddp_rd_overw), .B1(yadd_b[6]));
oai221x2_hvt I86_1_ ( .C0(yadd_b[8]), .A1(net565), .Y(yp1_sel_b[1]),
     .A0(yadd_b[7]), .B0(vddp_rd_overw), .B1(yadd[6]));
oai221x2_hvt I86_0_ ( .C0(yadd_b[8]), .A1(net565), .Y(yp1_sel_b[0]),
     .A0(yadd_b[7]), .B0(vddp_rd_overw), .B1(yadd_b[6]));
vdd_tiehigh I198 ( .vdd_tieh(vdd_tieh));
exor2_hvt I151_3_ ( .A(net339[0]), .Y(sb25low_b[3]), .B(pgm_hvact_b));
exor2_hvt I151_2_ ( .A(net339[1]), .Y(sb25low_b[2]), .B(pgm_hvact_b));
exor2_hvt I151_1_ ( .A(net339[2]), .Y(sb25low_b[1]), .B(pgm_hvact_b));
exor2_hvt I151_0_ ( .A(net339[3]), .Y(sb25low_b[0]), .B(pgm_hvact_b));
anor21_hvt I119_1_ ( .A(fsm_rowadd[1]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I119_0_ ( .A(fsm_rowadd[0]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
anor21_hvt I109 ( .A(pgm_hvact), .B(fsm_tm_allwl_h), .Y(net394),
     .C(nvcmen_buf_b));
ml_ls_vdd2vdd25 I168_3_ ( .in(net411[0]), .sup(vddp_),
     .out_vddio_b(sb25_high_25[3]), .out_vddio(net299[0]),
     .in_b(net552[0]));
ml_ls_vdd2vdd25 I168_2_ ( .in(net411[1]), .sup(vddp_),
     .out_vddio_b(sb25_high_25[2]), .out_vddio(net299[1]),
     .in_b(net552[1]));
ml_ls_vdd2vdd25 I168_1_ ( .in(net411[2]), .sup(vddp_),
     .out_vddio_b(sb25_high_25[1]), .out_vddio(net299[2]),
     .in_b(net552[2]));
ml_ls_vdd2vdd25 I168_0_ ( .in(net411[3]), .sup(vddp_),
     .out_vddio_b(sb25_high_25[0]), .out_vddio(net299[3]),
     .in_b(net552[3]));
ml_ls_vdd2vdd25 I167_3_ ( .in(net407[0]), .sup(vddp_),
     .out_vddio_b(sb25_gnd_25[3]), .out_vddio(net304[0]),
     .in_b(net549[0]));
ml_ls_vdd2vdd25 I167_2_ ( .in(net407[1]), .sup(vddp_),
     .out_vddio_b(sb25_gnd_25[2]), .out_vddio(net304[1]),
     .in_b(net549[1]));
ml_ls_vdd2vdd25 I167_1_ ( .in(net407[2]), .sup(vddp_),
     .out_vddio_b(sb25_gnd_25[1]), .out_vddio(net304[2]),
     .in_b(net549[2]));
ml_ls_vdd2vdd25 I167_0_ ( .in(net407[3]), .sup(vddp_),
     .out_vddio_b(sb25_gnd_25[0]), .out_vddio(net304[3]),
     .in_b(net549[3]));
ml_ls_vdd2vdd25 I144_3_ ( .in(net387[0]), .sup(vddp_),
     .out_vddio_b(sbhv_high_25[3]), .out_vddio(net522[0]),
     .in_b(net544[0]));
ml_ls_vdd2vdd25 I144_2_ ( .in(net387[1]), .sup(vddp_),
     .out_vddio_b(sbhv_high_25[2]), .out_vddio(net522[1]),
     .in_b(net544[1]));
ml_ls_vdd2vdd25 I144_1_ ( .in(net387[2]), .sup(vddp_),
     .out_vddio_b(sbhv_high_25[1]), .out_vddio(net522[2]),
     .in_b(net544[2]));
ml_ls_vdd2vdd25 I144_0_ ( .in(net387[3]), .sup(vddp_),
     .out_vddio_b(sbhv_high_25[0]), .out_vddio(net522[3]),
     .in_b(net544[3]));
ml_ls_vdd2vdd25 I148_3_ ( .in(net393[0]), .sup(vddp_),
     .out_vddio_b(sbhv_gnd_25[3]), .out_vddio(net523[0]),
     .in_b(net546[0]));
ml_ls_vdd2vdd25 I148_2_ ( .in(net393[1]), .sup(vddp_),
     .out_vddio_b(sbhv_gnd_25[2]), .out_vddio(net523[1]),
     .in_b(net546[1]));
ml_ls_vdd2vdd25 I148_1_ ( .in(net393[2]), .sup(vddp_),
     .out_vddio_b(sbhv_gnd_25[1]), .out_vddio(net523[2]),
     .in_b(net546[2]));
ml_ls_vdd2vdd25 I148_0_ ( .in(net393[3]), .sup(vddp_),
     .out_vddio_b(sbhv_gnd_25[0]), .out_vddio(net523[3]),
     .in_b(net546[3]));
ml_pump_a_clkdly I141_3_ ( .in(net393[0]), .out(net317[0]));
ml_pump_a_clkdly I141_2_ ( .in(net393[1]), .out(net317[1]));
ml_pump_a_clkdly I141_1_ ( .in(net393[2]), .out(net317[2]));
ml_pump_a_clkdly I141_0_ ( .in(net393[3]), .out(net317[3]));
ml_pump_a_clkdly I219_3_ ( .in(net387[0]), .out(net319[0]));
ml_pump_a_clkdly I219_2_ ( .in(net387[1]), .out(net319[1]));
ml_pump_a_clkdly I219_1_ ( .in(net387[2]), .out(net319[2]));
ml_pump_a_clkdly I219_0_ ( .in(net387[3]), .out(net319[3]));
ml_pump_a_clkdly I169_3_ ( .in(net411[0]), .out(net321[0]));
ml_pump_a_clkdly I169_2_ ( .in(net411[1]), .out(net321[1]));
ml_pump_a_clkdly I169_1_ ( .in(net411[2]), .out(net321[2]));
ml_pump_a_clkdly I169_0_ ( .in(net411[3]), .out(net321[3]));
ml_pump_a_clkdly I170_3_ ( .in(net407[0]), .out(net323[0]));
ml_pump_a_clkdly I170_2_ ( .in(net407[1]), .out(net323[1]));
ml_pump_a_clkdly I170_1_ ( .in(net407[2]), .out(net323[2]));
ml_pump_a_clkdly I170_0_ ( .in(net407[3]), .out(net323[3]));
nor3_hvt I111 ( .B(fsm_tm_allbl_l), .Y(yp3_b_high_b),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_l));
nor3_hvt I112 ( .C(yp3_b_high_b), .A(nvcmen_buf_b), .B(fsm_tm_allbl_h),
     .Y(net331));
nor3_hvt I57 ( .C(fsm_tm_allbl_h), .A(fsm_tm_allbl_l),
     .B(fsm_tm_testdec), .Y(net335));
anor31_hvt I155_3_ ( .A(ensb25_dec), .D(net395), .B(xadd[1]),
     .Y(net339[0]), .C(xadd[0]));
anor31_hvt I155_2_ ( .A(ensb25_dec), .D(net395), .B(xadd[1]),
     .Y(net339[1]), .C(xadd_b[0]));
anor31_hvt I155_1_ ( .A(ensb25_dec), .D(net395), .B(xadd_b[1]),
     .Y(net339[2]), .C(xadd[0]));
anor31_hvt I155_0_ ( .A(ensb25_dec), .D(net395), .B(xadd_b[1]),
     .Y(net339[3]), .C(xadd_b[0]));
anor31_hvt I121_3_ ( .A(net397), .D(net399), .B(xadd[1]),
     .Y(sbhvlow_b[3]), .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net397), .D(net399), .B(xadd[1]),
     .Y(sbhvlow_b[2]), .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net397), .D(net399), .B(xadd_b[1]),
     .Y(sbhvlow_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net397), .D(net399), .B(xadd_b[1]),
     .Y(sbhvlow_b[0]), .C(xadd_b[0]));
anor31_hvt I107 ( .A(fsm_tm_testdec), .D(net331), .B(nvcmen_buf),
     .Y(net349), .C(yadd[0]));
anor31_hvt I108 ( .A(fsm_tm_testdec), .D(net331), .B(nvcmen_buf),
     .Y(net354), .C(yadd_b[0]));
oai22x2_hvt I93 ( .A1(net381), .Y(net357), .A0(net453),
     .B0(fsm_nv_rri_trim), .B1(fsm_nv_sisi_ui));
nand4_hvt I122 ( .D(fsm_lshven), .C(pgm_hvact), .A(tm_allwl_l_b),
     .Y(net396), .B(blk_dec));
nand4_hvt I49_7_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[7]), .B(yadd[2]));
nand4_hvt I49_6_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[6]), .B(yadd[2]));
nand4_hvt I49_5_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[5]), .B(yadd[2]));
nand4_hvt I49_4_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[4]), .B(yadd[2]));
nand4_hvt I49_3_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[3]), .B(yadd_b[2]));
nand4_hvt I49_2_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[2]), .B(yadd_b[2]));
nand4_hvt I49_1_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[1]), .B(yadd_b[2]));
nand4_hvt I49_0_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[0]), .B(yadd_b[2]));
nand4_hvt I27 ( .D(fsm_blkadd[0]), .Y(blk_dec_b), .B(fsm_blkadd[2]),
     .C(fsm_blkadd[1]), .A(fsm_blkadd[3]));
inv_hvt I207 ( .A(net0579), .Y(ref_pgm));
inv_hvt I200 ( .A(fsm_tm_testdec), .Y(net377));
inv_hvt I120_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I120_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I181 ( .A(all_blk_sel_b), .Y(net381));
inv_hvt I161 ( .A(net570), .Y(net383));
inv_hvt I158 ( .A(pgm_hvact_b), .Y(pgm_hvact));
inv_hvt I142_3_ ( .A(net544[0]), .Y(net387[0]));
inv_hvt I142_2_ ( .A(net544[1]), .Y(net387[1]));
inv_hvt I142_1_ ( .A(net544[2]), .Y(net387[2]));
inv_hvt I142_0_ ( .A(net544[3]), .Y(net387[3]));
inv_hvt I157 ( .A(fsm_pgmvfy), .Y(net389));
inv_hvt I134_3_ ( .A(sbhvlow_b[3]), .Y(net391[0]));
inv_hvt I134_2_ ( .A(sbhvlow_b[2]), .Y(net391[1]));
inv_hvt I134_1_ ( .A(sbhvlow_b[1]), .Y(net391[2]));
inv_hvt I134_0_ ( .A(sbhvlow_b[0]), .Y(net391[3]));
inv_hvt I143_3_ ( .A(net546[0]), .Y(net393[0]));
inv_hvt I143_2_ ( .A(net546[1]), .Y(net393[1]));
inv_hvt I143_1_ ( .A(net546[2]), .Y(net393[2]));
inv_hvt I143_0_ ( .A(net546[3]), .Y(net393[3]));
inv_hvt I160 ( .A(net394), .Y(net395));
inv_hvt I123 ( .A(net396), .Y(net397));
inv_hvt I125 ( .A(net490), .Y(net399));
inv_hvt I189 ( .A(fsm_nvcmen), .Y(nvcmen_buf_b));
inv_hvt I164 ( .A(net402), .Y(net403));
inv_hvt I131 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I171_3_ ( .A(net549[0]), .Y(net407[0]));
inv_hvt I171_2_ ( .A(net549[1]), .Y(net407[1]));
inv_hvt I171_1_ ( .A(net549[2]), .Y(net407[2]));
inv_hvt I171_0_ ( .A(net549[3]), .Y(net407[3]));
inv_hvt I172_3_ ( .A(sb25low_b[3]), .Y(net409[0]));
inv_hvt I172_2_ ( .A(sb25low_b[2]), .Y(net409[1]));
inv_hvt I172_1_ ( .A(sb25low_b[1]), .Y(net409[2]));
inv_hvt I172_0_ ( .A(sb25low_b[0]), .Y(net409[3]));
inv_hvt I173_3_ ( .A(net552[0]), .Y(net411[0]));
inv_hvt I173_2_ ( .A(net552[1]), .Y(net411[1]));
inv_hvt I173_1_ ( .A(net552[2]), .Y(net411[2]));
inv_hvt I173_0_ ( .A(net552[3]), .Y(net411[3]));
inv_hvt I97 ( .A(fsm_multibl_read), .Y(net413));
inv_hvt I94 ( .A(net357), .Y(vddp_rd_overw));
inv_hvt I84 ( .A(nvcmen_buf_b), .Y(nvcmen_buf));
inv_hvt I72_7_ ( .A(yp2_sel_b[7]), .Y(yp2_sel[7]));
inv_hvt I72_6_ ( .A(yp2_sel_b[6]), .Y(yp2_sel[6]));
inv_hvt I72_5_ ( .A(yp2_sel_b[5]), .Y(yp2_sel[5]));
inv_hvt I72_4_ ( .A(yp2_sel_b[4]), .Y(yp2_sel[4]));
inv_hvt I72_3_ ( .A(yp2_sel_b[3]), .Y(yp2_sel[3]));
inv_hvt I72_2_ ( .A(yp2_sel_b[2]), .Y(yp2_sel[2]));
inv_hvt I72_1_ ( .A(yp2_sel_b[1]), .Y(yp2_sel[1]));
inv_hvt I72_0_ ( .A(yp2_sel_b[0]), .Y(yp2_sel[0]));
inv_hvt I66 ( .A(net349), .Y(net622));
inv_hvt I46_8_ ( .A(fsm_coladd[8]), .Y(yadd_b[8]));
inv_hvt I46_7_ ( .A(fsm_coladd[7]), .Y(yadd_b[7]));
inv_hvt I46_6_ ( .A(fsm_coladd[6]), .Y(yadd_b[6]));
inv_hvt I46_5_ ( .A(fsm_coladd[5]), .Y(yadd_b[5]));
inv_hvt I46_4_ ( .A(fsm_coladd[4]), .Y(yadd_b[4]));
inv_hvt I46_3_ ( .A(fsm_coladd[3]), .Y(yadd_b[3]));
inv_hvt I46_2_ ( .A(fsm_coladd[2]), .Y(yadd_b[2]));
inv_hvt I46_1_ ( .A(fsm_coladd[1]), .Y(yadd_b[1]));
inv_hvt I46_0_ ( .A(fsm_coladd[0]), .Y(yadd_b[0]));
inv_hvt I201 ( .A(fsm_tm_rd_mode), .Y(net425));
inv_hvt I25_2_ ( .A(tdec_b[2]), .Y(tdec[2]));
inv_hvt I25_1_ ( .A(tdec_b[1]), .Y(tdec[1]));
inv_hvt I25_0_ ( .A(tdec_b[0]), .Y(tdec[0]));
inv_hvt I24_2_ ( .A(net629[0]), .Y(tdec_b[2]));
inv_hvt I24_1_ ( .A(net629[1]), .Y(tdec_b[1]));
inv_hvt I24_0_ ( .A(net629[2]), .Y(tdec_b[0]));
inv_hvt I38_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I38_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I38_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I40 ( .A(net591), .Y(sa_bl_to_pgm_glb));
inv_hvt I103 ( .A(net511), .Y(en_blinhi_pgm_b));
inv_hvt I47_8_ ( .A(yadd_b[8]), .Y(yadd[8]));
inv_hvt I47_7_ ( .A(yadd_b[7]), .Y(yadd[7]));
inv_hvt I47_6_ ( .A(yadd_b[6]), .Y(yadd[6]));
inv_hvt I47_5_ ( .A(yadd_b[5]), .Y(yadd[5]));
inv_hvt I47_4_ ( .A(yadd_b[4]), .Y(yadd[4]));
inv_hvt I47_3_ ( .A(yadd_b[3]), .Y(yadd[3]));
inv_hvt I47_2_ ( .A(yadd_b[2]), .Y(yadd[2]));
inv_hvt I47_1_ ( .A(yadd_b[1]), .Y(yadd[1]));
inv_hvt I47_0_ ( .A(yadd_b[0]), .Y(yadd[0]));
inv_hvt I71 ( .A(net500), .Y(yp21_b_low_b));
inv_hvt I51_7_ ( .A(yp3_sel_b[7]), .Y(yp3_sel[7]));
inv_hvt I51_6_ ( .A(yp3_sel_b[6]), .Y(yp3_sel[6]));
inv_hvt I51_5_ ( .A(yp3_sel_b[5]), .Y(yp3_sel[5]));
inv_hvt I51_4_ ( .A(yp3_sel_b[4]), .Y(yp3_sel[4]));
inv_hvt I51_3_ ( .A(yp3_sel_b[3]), .Y(yp3_sel[3]));
inv_hvt I51_2_ ( .A(yp3_sel_b[2]), .Y(yp3_sel[2]));
inv_hvt I51_1_ ( .A(yp3_sel_b[1]), .Y(yp3_sel[1]));
inv_hvt I51_0_ ( .A(yp3_sel_b[0]), .Y(yp3_sel[0]));
inv_hvt I61 ( .A(net594), .Y(net443));
inv_hvt I28 ( .A(blk_dec_b), .Y(blk_dec));
inv_hvt I69 ( .A(net354), .Y(net612));
inv_hvt I117_1_ ( .A(yp_test_b[1]), .Y(yp_test[1]));
inv_hvt I117_0_ ( .A(yp_test_b[0]), .Y(yp_test[0]));
inv_hvt I185 ( .A(tm_tcol), .Y(net451));
inv_hvt I90 ( .A(net562), .Y(net453));
inv_25 I104 ( .IN(net606), .OUT(en_blinhi_pgm_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net620), .OUT(yp3_b_high_even_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I79 ( .IN(net610), .OUT(yp3_b_high_odd_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I77 ( .IN(net615), .OUT(yp3_b_low_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
nand3_hvt I204 ( .Y(yp1_sel_b[4]), .B(yadd_b[7]), .C(yadd[8]),
     .A(yadd_b[6]));
nand3_hvt I205 ( .Y(yp1_sel_b[5]), .B(yadd_b[7]), .C(yadd[6]),
     .A(yadd[8]));
nand3_hvt I156 ( .Y(pgm_hvact_b), .B(fsm_pgm), .C(net389),
     .A(fsm_lshven));
nand3_hvt I127 ( .Y(net490), .B(pgm_hvact), .C(fsm_tm_allwl_h),
     .A(fsm_lshven));
nand3_hvt I163 ( .C(tm_allwl_l_b), .A(fsm_vpxaset), .Y(net402),
     .B(sa_bl_to_blsa));
nand3_hvt I70 ( .C(nvcmen_buf), .A(net588), .Y(net500), .B(net377));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(tdec[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(tdec[1]), .C(tdec_b[0]),
     .A(tdec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(tdec_b[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I73_7_ ( .A(yadd[5]), .C(yadd[3]), .Y(yp2_sel_b[7]),
     .B(yadd[4]));
nand3_hvt I73_6_ ( .A(yadd[5]), .C(yadd_b[3]), .Y(yp2_sel_b[6]),
     .B(yadd[4]));
nand3_hvt I73_5_ ( .A(yadd[5]), .C(yadd[3]), .Y(yp2_sel_b[5]),
     .B(yadd_b[4]));
nand3_hvt I73_4_ ( .A(yadd[5]), .C(yadd_b[3]), .Y(yp2_sel_b[4]),
     .B(yadd_b[4]));
nand3_hvt I73_3_ ( .A(yadd_b[5]), .C(yadd[3]), .Y(yp2_sel_b[3]),
     .B(yadd[4]));
nand3_hvt I73_2_ ( .A(yadd_b[5]), .C(yadd_b[3]), .Y(yp2_sel_b[2]),
     .B(yadd[4]));
nand3_hvt I73_1_ ( .A(yadd_b[5]), .C(yadd[3]), .Y(yp2_sel_b[1]),
     .B(yadd_b[4]));
nand3_hvt I73_0_ ( .A(yadd_b[5]), .C(yadd_b[3]), .Y(yp2_sel_b[0]),
     .B(yadd_b[4]));
nor4_hvt I98 ( .B(fsm_tm_allbl_l), .Y(net511), .D(nvcmen_buf_b),
     .A(net573), .C(fsm_tm_allbl_l));
nor4_hvt I52 ( .D(net580), .B(fsm_tm_allbl_h), .Y(ymux_dis_b),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_h));
nor2_hvt I202 ( .A(yp1_sel_b[4]), .B(tm_tcol), .Y(yp1_sel[4]));
nor2_hvt I203 ( .A(yp1_sel_b[5]), .B(tm_tcol), .Y(yp1_sel[5]));
nor2_hvt I195 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I128_3_ ( .B(net317[0]), .A(net391[0]), .Y(net544[0]));
nor2_hvt I128_2_ ( .B(net317[1]), .A(net391[1]), .Y(net544[1]));
nor2_hvt I128_1_ ( .B(net317[2]), .A(net391[2]), .Y(net544[2]));
nor2_hvt I128_0_ ( .B(net317[3]), .A(net391[3]), .Y(net544[3]));
nor2_hvt I140_3_ ( .A(net319[0]), .Y(net546[0]), .B(sbhvlow_b[3]));
nor2_hvt I140_2_ ( .A(net319[1]), .Y(net546[1]), .B(sbhvlow_b[2]));
nor2_hvt I140_1_ ( .A(net319[2]), .Y(net546[2]), .B(sbhvlow_b[1]));
nor2_hvt I140_0_ ( .A(net319[3]), .Y(net546[3]), .B(sbhvlow_b[0]));
nor2_hvt I176_3_ ( .A(sb25low_b[3]), .Y(net549[0]), .B(net321[0]));
nor2_hvt I176_2_ ( .A(sb25low_b[2]), .Y(net549[1]), .B(net321[1]));
nor2_hvt I176_1_ ( .A(sb25low_b[1]), .Y(net549[2]), .B(net321[2]));
nor2_hvt I176_0_ ( .A(sb25low_b[0]), .Y(net549[3]), .B(net321[3]));
nor2_hvt I177_3_ ( .A(net323[0]), .Y(net552[0]), .B(net409[0]));
nor2_hvt I177_2_ ( .A(net323[1]), .Y(net552[1]), .B(net409[1]));
nor2_hvt I177_1_ ( .A(net323[2]), .Y(net552[2]), .B(net409[2]));
nor2_hvt I177_0_ ( .A(net323[3]), .Y(net552[3]), .B(net409[3]));
nor2_hvt I114 ( .A(tm_tcol), .B(net600), .Y(ymux_en_core));
nor2_hvt I186 ( .A(net451), .B(net600), .Y(ymux_test_en));
nor2_hvt I88 ( .A(fsm_tm_rd_mode), .B(fsm_pgmvfy), .Y(net562));
nor2_hvt I96 ( .A(net357), .B(net413), .Y(net565));
nor2_hvt I75_3_ ( .A(yp1_sel_b[3]), .B(tm_tcol), .Y(yp1_sel[3]));
nor2_hvt I75_2_ ( .A(yp1_sel_b[2]), .B(tm_tcol), .Y(yp1_sel[2]));
nor2_hvt I75_1_ ( .A(yp1_sel_b[1]), .B(tm_tcol), .Y(yp1_sel[1]));
nor2_hvt I75_0_ ( .A(yp1_sel_b[0]), .B(tm_tcol), .Y(yp1_sel[0]));
nor2_hvt I206 ( .A(fsm_pgmvfy), .B(fsm_pgm), .Y(net0579));
nand2_hvt I162 ( .A(blk_dec), .Y(net570), .B(tm_allwl_l_b));
nand2_hvt I101 ( .A(pgm_hvact), .Y(net573), .B(pgm_hvact));
nand2_hvt I35 ( .B(one_blk_sel_b), .Y(sa_bl_to_blsa),
     .A(all_blk_sel_b));
nand2_hvt I53 ( .A(fsm_nvcmen), .B(fsm_lshven), .Y(net580));
nand2_hvt I116_1_ ( .A(yadd[0]), .Y(yp_test_b[1]), .B(ymux_test_en));
nand2_hvt I116_0_ ( .A(yadd_b[0]), .Y(yp_test_b[0]), .B(ymux_test_en));
nand2_hvt I59 ( .A(fsm_lshven), .Y(net588), .B(pgm_hvact));
nand2_hvt I39 ( .A(blk_dec), .Y(net591), .B(fsm_pgmien));
nand2_hvt I60 ( .A(net588), .Y(net594), .B(net335));
nand2_hvt I89 ( .A(fsm_tm_rd_mode), .Y(one_blk_sel_b), .B(blk_dec));
oai21x2_hvt I55 ( .A1(sa_bl_to_blsa), .Y(net600), .A0(blk_dec),
     .B0(ymux_dis_b));
ml_ls_vdd25_nor2 I106 ( .in(net511), .sup(ysup_25),
     .out_vddio_b(net605), .out_vddio(net606), .in_b(en_blinhi_pgm_b));
ml_ls_vdd25_nor2 I68 ( .in(net354), .sup(ysup_25),
     .out_vddio_b(net610), .out_vddio(net611), .in_b(net612));
ml_ls_vdd25_nor2 I192 ( .in(net594), .sup(ysup_25),
     .out_vddio_b(net615), .out_vddio(net616), .in_b(net443));
ml_ls_vdd25_nor2 I65 ( .in(net349), .sup(ysup_25),
     .out_vddio_b(net620), .out_vddio(net621), .in_b(net622));
mux2_hvt I152 ( .in1(net383), .in0(net403), .out(ensb25_dec),
     .sel(pgm_hvact));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net629[0]), .sel(ref_pgm));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net629[1]), .sel(ref_pgm));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net629[2]), .sel(ref_pgm));

endmodule
// Library - NVCM, Cell - ml_core_sa_resbot_m2, View - schematic
// LAST TIME SAVED: Sep 11 10:45:00 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa_resbot_m2 ( bl_in, bl_out, div_2r, div_3r, nwell,
     sa_ngate_25, sa_pgate_vpxa );
inout  bl_in, bl_out, div_2r, div_3r, nwell;


input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M4 ( .D(net115), .B(gnd_), .G(sa_ngate_25[4]), .S(bl_out));
nch_25  M3 ( .D(net090), .B(gnd_), .G(sa_ngate_25[3]), .S(net115));
nch_25  M0 ( .D(net086), .B(gnd_), .G(sa_ngate_25[2]), .S(net090));
nch_25  M32 ( .D(net111), .B(gnd_), .G(sa_ngate_25[1]), .S(net086));
pch_25  M5 ( .D(bl_out), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net115));
pch_25  M1 ( .D(net090), .B(nwell), .G(sa_pgate_vpxa[2]), .S(net086));
pch_25  M2 ( .D(net115), .B(nwell), .G(sa_pgate_vpxa[3]), .S(net090));
pch_25  M37 ( .D(net086), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net111));
rppolywo_m  R31 ( .MINUS(net099), .PLUS(div_3r), .BULK(gnd_));
rppolywo_m  R32 ( .MINUS(div_2r), .PLUS(net099), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(div_3r), .PLUS(net111), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net111), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R30 ( .MINUS(net0111), .PLUS(div_2r), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(bl_out), .PLUS(net0111), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa_refres, View - schematic
// LAST TIME SAVED: Sep 11 10:40:27 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa_refres ( bot, nwell, wp_ref, sa_ngate_25,
     sa_pgate_vpxa );
inout  bot, nwell, wp_ref;


input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M32 ( .D(net44), .B(gnd_), .G(sa_ngate_25[1]), .S(net40));
nch_25  M2 ( .D(net50), .B(gnd_), .G(sa_ngate_25[3]), .S(net084));
nch_25  M6 ( .D(net084), .B(gnd_), .G(sa_ngate_25[4]), .S(bot));
nch_25  M1 ( .D(net40), .B(gnd_), .G(sa_ngate_25[2]), .S(net50));
pch_25  M3 ( .D(net084), .B(nwell), .G(sa_pgate_vpxa[3]), .S(net50));
pch_25  M37 ( .D(net40), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net44));
pch_25  M5 ( .D(bot), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net084));
pch_25  M0 ( .D(net50), .B(nwell), .G(sa_pgate_vpxa[2]), .S(net40));
rppolywo_m  R2 ( .MINUS(net096), .PLUS(net090), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(bot), .PLUS(net32), .BULK(gnd_));
rppolywo_m  R6 ( .MINUS(net32), .PLUS(net096), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net090), .PLUS(net44), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net44), .PLUS(wp_ref), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa_resbot, View - schematic
// LAST TIME SAVED: Apr  9 15:18:14 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa_resbot ( bl_in, bl_out, div_2r, div_3r, nwell,
     sa_ngate_25, sa_pgate_vpxa );
inout  bl_in, bl_out, div_2r, div_3r, nwell;


input [4:1]  sa_pgate_vpxa;
input [4:1]  sa_ngate_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M4 ( .D(net115), .B(gnd_), .G(sa_ngate_25[4]), .S(bl_out));
nch_25  M3 ( .D(div_2r), .B(gnd_), .G(sa_ngate_25[3]), .S(net115));
nch_25  M0 ( .D(div_3r), .B(gnd_), .G(sa_ngate_25[2]), .S(div_2r));
nch_25  M32 ( .D(net111), .B(gnd_), .G(sa_ngate_25[1]), .S(div_3r));
pch_25  M5 ( .D(bl_out), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net115));
pch_25  M1 ( .D(div_2r), .B(nwell), .G(sa_pgate_vpxa[2]), .S(div_3r));
pch_25  M2 ( .D(net115), .B(nwell), .G(sa_pgate_vpxa[3]), .S(div_2r));
pch_25  M37 ( .D(div_3r), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net111));
rppolywo_m  R31 ( .MINUS(net099), .PLUS(div_3r), .BULK(gnd_));
rppolywo_m  R32 ( .MINUS(div_2r), .PLUS(net099), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(div_3r), .PLUS(net111), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net111), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R30 ( .MINUS(net115), .PLUS(div_2r), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(bl_out), .PLUS(net115), .BULK(gnd_));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Aug  3 14:03:13 2007
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module sbtlibn65lp_ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp, View - schematic
// LAST TIME SAVED: Jan 21 17:21:12 2008
// NETLIST TIME: Aug 24 09:58:58 2009
`timescale 1ns / 1ns 

module ml_core_sa_comp ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_b_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M4_1_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M0 ( .D(out_div), .B(vddp_), .G(in_div), .S(net65));
pch_25  M3 ( .D(out_ref), .B(vddp_), .G(in_ref), .S(net65));
nch_25  M1 ( .D(out_ref), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M2 ( .D(out_div), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M8 ( .D(out_ref), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M5 ( .D(out_div), .B(GND_), .G(saen_b_25), .S(gnd_));

endmodule
// Library - io, Cell - PDT08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 15:32:26 2007
// NETLIST TIME: Aug 24 09:58:57 2009
`timescale 1ns / 1ns 

module PDT08DGZ ( PAD, I, OEN );
inout  PAD;

input  I, OEN;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
