---------------------------------------------------------------------------
---------------------------------------------------------------------------
--
--      IO LOGIC MODULE
--
--      FOR IPRO INDUSTRIAL FPGA
--
--      VHDL DESIGN FILE :IOLOGIC10.VHD
--
--      by: M. Stamer
--      VIDEOJET TECHNOLOGIES INC.
--
---------------------------------------------------------------------------
---------------------------------------------------------------------------
--
-------------------------------------------------------------------------------
--
-- Copyright 2002 Videojet Technologies Inc. All Rights Reserved. 
--
-- An unpublished work of Videojet Technologies Inc. The software and 
-- documentation contained herein are copyrighted works which include 
-- confidential information and trade secrets proprietary to Videojet 
-- Technologies Inc. and shall not be copied, duplicated, disclosed or used, 
-- in whole or in part, except pursuant to the License Agreement or as 
-- otherwise expressly approved by Videojet Technologies Inc.
--
-------------------------------------------------------------------------------
-- This module implements the I/O functions for the revised IPRO-2
-- printer.  In this design, each of the general purpose inputs
-- has software configurable function and assignment.  Inputs can
-- be configured for polarity, one of four choices of digital filtering
-- or grouped for any change (after debounce/filtering) to cause an
-- interrupt.
--
-- Each general purpose output is also configurable to be generated by
-- a software selected function.  Output polarity is always active low.
--
-- All configuring of inputs and outputs is done by means of software
-- writing to configuration registers.

-- Modified for use with Synplicity synthesis software.

-- IOLOGIC3.VHD modified to support selective interrupt clear and
-- flag clear.  This was implemented by gating the respective clear
-- command with the appropriate data bit for each input interrupt
-- entity.  Also corrected input edge select to be always leading
-- edge for most inputs.  In addition, added prod3, which has an
-- additional input to enable generation of interrupts on both edges
-- of input.

-- IOLOGIC4.VHD revised (and simplified) the gated output control
-- logic options.

-- IOLOGIC5.VHD revised the pulsed output feature to trigger based on the
-- writing of ones at the specific bits and not requiring the writing of a
-- zero to enable the writing of a subsequent one to trigger the next pulse.

-- IOLOGIC6.VHD corrected the general input organization in realigning
-- which input corresponded to the opto-isolated inputs and thus, the
-- corresponding software gating features.

-- IOLOGIC7.VHD adds the abilitoy to re-trigger the one-shot timers prior to
-- the expiration of their timeout period. 
--
--  Also corrected the polarity of the gating signals for gated outputs and
--  corrected which outputs are gated.
--
-- IOLOGIC8.VHD was downsized for the Low-End CIJ printer.  
--
-- IOLOGIC9.VHD is an expanded version of IOLOGIC7.VHD.  This module is the
-- starting IO module for the Videojet 1000 printer (platform).  Here, the number of
-- inputs and outputs is expanded to match the new IO Expansion board.  IO
-- assumptions are similar to IPRO2, in lueue of any concrete FRS.  Known changes
-- include a single printhead, two PDs, 11 general inputs, 9 general outputs.
-- Whether or not a product uses these features will be determined under
-- software control.  A new input, not part of this module, senses the 
-- presence of an IO expansion board.  For now, the upper one or two inputs
-- will be used to indicate which type of IO module is attached.
-- 
-- This version of IOLOGIC9 (file called IOLOGIC_IPRO2.VHD), uses only the IPRO2 
-- level of IO functionality.  The other IO pins are used for:
	-- A. selection inputs for expansion board type;
	-- B. simple port control or duplication of other inputs or outputs; i.e.
	--    not customized parameters.
--	
-- The first attempt fitting result with this file allowed the total FPGA design
-- to just fit into an Altera ACEX1K30 size part, but using 1706 out of 1728 available
-- logic cells.  This still did not include the finalized KBD logic or expansion
-- board select pins ( a minor impact).  Thus, we could save several dollars in
-- board cost if we standardize on the smaller FPGA.  Then, if a deluxe version
-- is needed, a new assembly version must be generated.
--
-- IOLOGIC10.VHD is the finalized IO interface plan for the VJ1000 controller.  This
-- will support nine inputs (8 message select inputs, one general purpose input) and 
-- eight outputs.  Most of the hardware support will reside on an optional expansion
-- card.  Three of these outputs are relay devices.  The tri-color alert light 
-- and siren connector are also supported.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

ENTITY iologic10 IS
    PORT(mclk, Nwr, Nreset, input_config1_dcd,
        output_config2_dcd,	outsrc_config3_dcd, outctrl_config4_dcd,
        intr_in_clr_dcd, flag_in_clr_dcd,
		clk1mh_tick, clk2kh_tick, clk2_9kh_tick, clk1_45kh_tick,
        clk362hz_tick, clk181hz_tick, print_enable1,
        image_done1 : in std_logic;

        Ngenin : in std_logic_vector(8 downto 0);

        data : in std_logic_vector(31 downto 0);

        Ngen_out : out std_logic_vector(7 downto 0);
        Ntri_red, Ntri_yel, Ntri_grn, Nsiren : out std_logic;
        
        input_filtered : out std_logic_vector(8 downto 0);
        intr_input_reg : out std_logic_vector(8 downto 0);
        input_flag_reg : out std_logic_vector(8 downto 0) );

END iologic10;

ARCHITECTURE archiologic10 OF iologic10 IS

--	attribute syn_hier of archiologic9 : architecture is "remove";

	SIGNAL input_config1, output_config2, outsrc_config3
        : std_logic_vector(31 downto 0);
	SIGNAL input_data, in_invreg, genin,
        inputreg2, inputreg3 : std_logic_vector(8 downto 0);
	SIGNAL output_data : std_logic_vector(7 downto 0);
	SIGNAL clk_div1 : std_logic_vector(3 downto 0);
	SIGNAL inputreg1 : std_logic_vector(9 downto 0);
	
	SIGNAL src_config0, src_config1, src_config2, src_config3,
        src_config4, src_config5, src_config6, src_config7, src_config8
		: std_logic_vector(1 downto 0); 
		
	SIGNAL count25, fltr_count, gatemode_a, gatemode_b 
		: std_logic_vector(2 downto 0);
		

    SIGNAL in_filter_select0, in_filter_select1,
        in_filter_select2, in_filter_select3, in_filter_select4, in_filter_select5,
        in_filter_select6, in_filter_select7, in_filter_select8, in_filter_select9,
        in_filter_select10, alert_data_red, alert_data_yel, alert_data_grn,
		alert_data_siren, pulse_width_0, pulse_width_1, pulse_width_2, pulse_width_3,
		pulse_width_4, pulse_width_5, pulse_width_6, pulse_width_7, pulse_width_8,
        mod_src_config0, mod_src_config1, mod_src_config2, mod_src_config3,
        mod_src_config4, mod_src_config5, mod_src_config6, mod_src_config7, 
		mod_src_config8 : std_logic_vector(1 downto 0);
			   
	SIGNAL flash_count : std_logic_vector(5 downto 0);

	SIGNAL input_filtered0_temp, input_filtered4_temp,
	input_config1_regen, output_config2_regen, outsrc_config3_regen,
	outctrl_config4_regen, intr_in_clr_regen, flag_in_clr_regen,
	clk8ms_del, clk8ms_tick, high, low, filter_regen, fltr2_5ms_tick,
    tick25, fltr_5ms_tick, fltr_10ms_tick, fltr_20ms_tick,
    fltr5mstick, fltr10mstick, fltr20mstick, count25_del, fltr_5ms_del, 
	fltr_10ms_del, fltr_20ms_del, flash_1sec, flash_half_sec, output_active,
	qtr_sec_toggle, half_sec_toggle, gate_enable_A, gate_enable_B, 
	out_enable0, out_enable1, out_enable2, out_enable3, 
    out_enable4, out_enable5, out_enable6, out_enable7, out_enable8,

    clock_choice0, intr_in0_enable,
    intr_in0_clr, flag_in0_clr, set_in0_overlap_fault,
    set_in0_bounce_warning, intr_in0_flag, intr_in0, in0_filtered,
    in0_edge_tick, 

    clock_choice1, intr_in1_enable,
    intr_in1_clr, flag_in1_clr, set_in1_overlap_fault,
    set_in1_bounce_warning, intr_in1_flag, intr_in1, in1_filtered,
    in1_edge_tick,

    clock_choice2, intr_in2_enable,
    intr_in2_clr, flag_in2_clr, set_in2_overlap_fault,
    set_in2_bounce_warning, intr_in2_flag, intr_in2, in2_filtered,
    in2_edge_tick,

    clock_choice3, intr_in3_enable,
    intr_in3_clr, flag_in3_clr, set_in3_overlap_fault,
    set_in3_bounce_warning, intr_in3_flag, intr_in3, in3_filtered,
    in3_edge_tick,

    clock_choice4, intr_in4_enable,
    intr_in4_clr, flag_in4_clr, set_in4_overlap_fault,
    set_in4_bounce_warning, intr_in4_flag, intr_in4, in4_filtered,
    in4_edge_tick,

    clock_choice5, intr_in5_enable,
    intr_in5_clr, flag_in5_clr, set_in5_overlap_fault,
    set_in5_bounce_warning, intr_in5_flag, intr_in5, in5_filtered,
    in5_edge_tick,

    clock_choice6, intr_in6_enable,
    intr_in6_clr, flag_in6_clr, set_in6_overlap_fault,
    set_in6_bounce_warning, intr_in6_flag, intr_in6, in6_filtered,
    in6_edge_tick,

    clock_choice7, intr_in7_enable,
    intr_in7_clr, flag_in7_clr, set_in7_overlap_fault,
    set_in7_bounce_warning, intr_in7_flag, intr_in7, in7_filtered,
    in7_edge_tick,

    clock_choice8, intr_in8_enable,
    intr_in8_clr, flag_in8_clr, set_in8_overlap_fault,
    set_in8_bounce_warning, intr_in8_flag, intr_in8, in8_filtered,
    in8_edge_tick,

--    clock_choice9, intr_in9_enable,
--    intr_in9_clr, flag_in9_clr, set_in9_overlap_fault,
--    set_in9_bounce_warning, intr_in9_flag, intr_in9, in9_filtered,
--    in9_edge_tick, 

--    clock_choice10, intr_in10_enable,
--    intr_in10_clr, flag_in10_clr, set_in10_overlap_fault,
--    set_in10_bounce_warning, intr_in10_flag, intr_in10, in10_filtered,
--    in10_edge_tick, 

    pulse_choice0, pulse_choice1, pulse_choice2, pulse_choice3,
    pulse_choice4, pulse_choice5, pulse_choice6, pulse_choice7, pulse_choice8,
    edge_out0, edge_out1, edge_out2, edge_out3,
    edge_out4, edge_out5, edge_out6, edge_out7, edge_out8, 
	two_edge_enable1, two_edge_enable3, 
    enabletick0, enabletick1, enabletick2, enabletick3, 
    enabletick4, enabletick5, enabletick6, enabletick7, enabletick8,
    out_choice0, out_choice1, out_choice2, out_choice3,
    out_choice4, out_choice5, out_choice6, out_choice7, out_choice8,
    out_choice_tick0, out_choice_tick1, out_choice_tick2, out_choice_tick3,
    out_choice_tick4, out_choice_tick5, out_choice_tick6, out_choice_tick7, 
	out_choice_tick8,
    out_choice_del0, out_choice_del1, out_choice_del2, out_choice_del3,
    out_choice_del4, out_choice_del5, out_choice_del6, out_choice_del7, 
	out_choice_del8,
    level_out0, level_out1, level_out2, level_out3,
    level_out4, level_out5, level_out6, level_out7, level_out8,
    gen_out0, gen_out1, gen_out2, gen_out3,
    gen_out4, gen_out5, gen_out6, gen_out7, gen_out8,
	pulse_mode_0, pulse_mode_1, pulse_mode_2, pulse_mode_3,
	pulse_mode_4, pulse_mode_5, pulse_mode_6, pulse_mode_7, pulse_mode_8,
    pulse_out0, pulse_out1, pulse_out2, pulse_out3,
    pulse_out4, pulse_out5, pulse_out6, pulse_out7, pulse_out8, tri_red, 
	tri_yel, tri_grn, siren : std_logic;

COMPONENT prod2
    PORT(mclk, Nreset, pd, pd_inv, pd_lead_edge_sel, enc_tick_choice,
		enable_in, pd_intr_clr, pd_flag_clr : in std_logic;
		set_pd_overlap_fault, set_pd_bounce_warning,
		pd_int_flag, pd_intr, pd_filtered, pd_edge_tick : out std_logic);
END COMPONENT;

--COMPONENT prod3
--    PORT(mclk, Nreset, pd, pd_inv, pd_lead_edge_sel, two_edge_enable, enc_tick_choice,
--		enable_in, pd_intr_clr, pd_flag_clr : in std_logic;
--		pd_int_flag, pd_intr, pd_filtered, pd_edge_tick : out std_logic);
--END COMPONENT;

COMPONENT pulse_5 IS PORT(mclk, Nreset, clk_tick, pulse_in : in std_logic;
		pulse_out : out std_logic);
    END COMPONENT;

COMPONENT pulse_rt_1ms IS PORT(mclk, Nreset, clk16kh_tick, pulse_in : in std_logic;
		pulse_out : out std_logic);
END COMPONENT;

COMPONENT selector_2 IS PORT(mclk, Nreset, enable, 
        input0, input1, selector: in std_logic;
		sel_out : out std_logic);
END COMPONENT;

COMPONENT selector_4
    PORT(mclk, Nreset, enable, 
        input0, input1, input2, input3: in std_logic;
        selector :std_logic_vector(1 downto 0);
		sel_out : out std_logic);
END COMPONENT;

	
     BEGIN
	genin(0) <= not Ngenin(0);		
	genin(1) <= not Ngenin(1);		
	genin(2) <= not Ngenin(2);		
	genin(3) <= not Ngenin(3);		
	genin(4) <= not Ngenin(4);		
	genin(5) <= not Ngenin(5);		
	genin(6) <= not Ngenin(6);		
	genin(7) <= not Ngenin(7);		
	genin(8) <= not Ngenin(8);	
--	genin(9) <= not Ngenin(9);	
--	genin(10) <= not Ngenin(10);	
	
	high <= '1';
	low  <= '0';

------------------- DIGITAL FILTER TIME BASE ---------------------

-- The input filtering and output pulse width timing is derived
-- using timing pulses generated in this section.  Input debounce
-- times will be software configurable individually for each input.
-- Output pulse or level mode is selectable.  If pulse mode is
-- selected, a selectable pulse width is generated.

    tick25 <= count25_del AND not(count25(2));

	timing2_5ms: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        fltr2_5ms_tick <= '0';
        count25 <= "000";
		count25_del <= '0';
	elsif(rising_edge (mclk)) then
        if(clk2kh_tick='1') then
            if(count25="100") then
                count25<="000";
            else
        	    count25 <= count25 + 1;
    	    end if;
	    end if;
        count25_del <= count25(2);
        fltr2_5ms_tick <= tick25;
	end if;
    END process timing2_5ms;


	timing_filter1: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        fltr_count <= "000";
	elsif(rising_edge (mclk)) then
        if(fltr2_5ms_tick='1') then
            fltr_count <= fltr_count + 1;
	    end if;
	end if;
    END process timing_filter1;

    fltr5mstick <= fltr_5ms_del AND not(fltr_count(0));
    fltr10mstick <= fltr_10ms_del AND not(fltr_count(1));
    fltr20mstick <= fltr_20ms_del AND not(fltr_count(2));

	timing_filter2: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        fltr_5ms_tick  <= '0';
        fltr_10ms_tick <= '0';
        fltr_20ms_tick <= '0';
        fltr_5ms_del  <= '0';
        fltr_10ms_del <= '0';
        fltr_20ms_del <= '0';
	elsif(rising_edge (mclk)) then
        fltr_5ms_del  <= fltr_count(0);
        fltr_10ms_del <= fltr_count(1);
        fltr_20ms_del <= fltr_count(2);
        fltr_5ms_tick  <= fltr5mstick;
        fltr_10ms_tick <= fltr10mstick;
        fltr_20ms_tick <= fltr20mstick;
	end if;
    END process timing_filter2;

------------------ INPUT FILTER CLOCK CHOICE --------------------
-- Syncronous multiplexer, one of four input pulse intervals
-- are selected based on configuration bits.

    mux0: selector_4 port map(mclk, Nreset, high,
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select0, clock_choice0);

    mux1: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select1, clock_choice1);

    mux2: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select2, clock_choice2);

    mux3: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select3, clock_choice3);

    mux4: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select4, clock_choice4);

    mux5: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select5, clock_choice5);

    mux6: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select6, clock_choice6);

    mux7: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select7, clock_choice7);

    mux8: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
        in_filter_select8, clock_choice8);

--    mux9: selector_4 port map(mclk, Nreset, high, 
--        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
--        in_filter_select9, clock_choice9);

--    mux10: selector_4 port map(mclk, Nreset, high, 
--        clk1mh_tick, fltr2_5ms_tick, fltr_5ms_tick, fltr_10ms_tick,
--        in_filter_select10, clock_choice10);


---------------------- INPUT FILTERING --------------------------

--        intr_in_clr_regen <= intr_in_clr_dcd AND not(Nwr);
        
        intr_in0_clr <= data(0) AND intr_in_clr_dcd AND not(Nwr);
        intr_in1_clr <= data(1) AND intr_in_clr_dcd AND not(Nwr);
        intr_in2_clr <= data(2) AND intr_in_clr_dcd AND not(Nwr);
        intr_in3_clr <= data(3) AND intr_in_clr_dcd AND not(Nwr);
        intr_in4_clr <= data(4) AND intr_in_clr_dcd AND not(Nwr);
        intr_in5_clr <= data(5) AND intr_in_clr_dcd AND not(Nwr);
        intr_in6_clr <= data(6) AND intr_in_clr_dcd AND not(Nwr);
        intr_in7_clr <= data(7) AND intr_in_clr_dcd AND not(Nwr);
        intr_in8_clr <= data(8) AND intr_in_clr_dcd AND not(Nwr);
--        intr_in9_clr <= data(9) AND intr_in_clr_dcd AND not(Nwr);
--        intr_in10_clr <= data(10) AND intr_in_clr_dcd AND not(Nwr);

--        flag_in_clr_regen <= flag_in_clr_dcd AND not(Nwr);

        flag_in0_clr <= data(0) AND flag_in_clr_dcd AND not(Nwr);
        flag_in1_clr <= data(1) AND flag_in_clr_dcd AND not(Nwr);
        flag_in2_clr <= data(2) AND flag_in_clr_dcd AND not(Nwr);
        flag_in3_clr <= data(3) AND flag_in_clr_dcd AND not(Nwr);
        flag_in4_clr <= data(4) AND flag_in_clr_dcd AND not(Nwr);
        flag_in5_clr <= data(5) AND flag_in_clr_dcd AND not(Nwr);
        flag_in6_clr <= data(6) AND flag_in_clr_dcd AND not(Nwr);
        flag_in7_clr <= data(7) AND flag_in_clr_dcd AND not(Nwr);
        flag_in8_clr <= data(8) AND flag_in_clr_dcd AND not(Nwr);
--        flag_in9_clr <= data(9) AND flag_in_clr_dcd AND not(Nwr);
--        flag_in10_clr <= data(10) AND flag_in_clr_dcd AND not(Nwr);


-- Note that IN3 and IN1 use prod3 instead of prod2.  This is
-- because certain FRS features require an interrupt on both
-- lead and trailing edges of certain inputs, if certain
-- features are selected.  Specifically, this includes use of
-- an input to enable/inhibit printing.  At other times, the same
-- input will be a normal input which can cause an interrupt
-- only on the lead edge transitions.

     in0: prod2 PORT MAP(
          mclk, Nreset, genin(0), in_invreg(0), high,
          clock_choice0, intr_in0_enable, intr_in0_clr, flag_in0_clr,
          set_in0_overlap_fault, set_in0_bounce_warning,
          intr_in0_flag, intr_in0, in0_filtered, in0_edge_tick);

     in1: prod2 PORT MAP(
          mclk, Nreset, genin(1), in_invreg(1), high,
          clock_choice1, intr_in1_enable, intr_in1_clr, flag_in1_clr,
          set_in1_overlap_fault, set_in1_bounce_warning,
          intr_in1_flag, intr_in1, in1_filtered, in1_edge_tick);

     in2: prod2 PORT MAP(
          mclk, Nreset, genin(2), in_invreg(2), high,
          clock_choice2, intr_in2_enable, intr_in2_clr, flag_in2_clr,
          set_in2_overlap_fault, set_in2_bounce_warning,
          intr_in2_flag, intr_in2, in2_filtered, in2_edge_tick);

     in3: prod2 PORT MAP(
          mclk, Nreset, genin(3), in_invreg(3), high,
          clock_choice3, intr_in3_enable, intr_in3_clr, flag_in3_clr,
          set_in3_overlap_fault, set_in3_bounce_warning,
          intr_in3_flag, intr_in3, in3_filtered, in3_edge_tick);

     in4: prod2 PORT MAP(
          mclk, Nreset, genin(4), in_invreg(4), high,
          clock_choice4, intr_in4_enable, intr_in4_clr, flag_in4_clr,
          set_in4_overlap_fault, set_in4_bounce_warning,
          intr_in4_flag, intr_in4, in4_filtered, in4_edge_tick);

     in5: prod2 PORT MAP(
          mclk, Nreset, genin(5), in_invreg(5), high,
          clock_choice5, intr_in5_enable, intr_in5_clr, flag_in5_clr,
          set_in5_overlap_fault, set_in5_bounce_warning,
          intr_in5_flag, intr_in5, in5_filtered, in5_edge_tick);

     in6: prod2 PORT MAP(
          mclk, Nreset, genin(6), in_invreg(6), high,
          clock_choice6, intr_in6_enable, intr_in6_clr, flag_in6_clr,
          set_in6_overlap_fault, set_in6_bounce_warning,
          intr_in6_flag, intr_in6, in6_filtered, in6_edge_tick);

     in7: prod2 PORT MAP(
          mclk, Nreset, genin(7), in_invreg(7), high, -- low,
          clock_choice7, intr_in7_enable, intr_in7_clr, flag_in7_clr,
          set_in7_overlap_fault, set_in7_bounce_warning,
          intr_in7_flag, intr_in7, in7_filtered, in7_edge_tick);

     in8: prod2 PORT MAP(
          mclk, Nreset, genin(8), in_invreg(8), high,
          clock_choice8, intr_in8_enable, intr_in8_clr, flag_in8_clr,
          set_in8_overlap_fault, set_in8_bounce_warning,
          intr_in8_flag, intr_in8, in8_filtered, in8_edge_tick);

--     in9: prod2 PORT MAP(
--          mclk, Nreset, genin(9), in_invreg(9), high, -- low,
--          clock_choice9, intr_in9_enable, intr_in9_clr, flag_in9_clr,
--          set_in9_overlap_fault, set_in9_bounce_warning,
--          intr_in9_flag, intr_in9, in9_filtered, in9_edge_tick);

--     in10: prod2 PORT MAP(
--          mclk, Nreset, genin(10), in_invreg(9), high, -- low,
--          clock_choice10, intr_in10_enable, intr_in10_clr, flag_in10_clr,
--          set_in10_overlap_fault, set_in10_bounce_warning,
--          intr_in10_flag, intr_in10, in10_filtered, in10_edge_tick);

          input_filtered0_temp <= in0_filtered;
          input_filtered(1) <= in1_filtered;
          input_filtered(2) <= in2_filtered;
          input_filtered(3) <= in3_filtered;
          input_filtered4_temp <= in4_filtered;
          input_filtered(5) <= in5_filtered;
          input_filtered(6) <= in6_filtered;
          input_filtered(7) <= in7_filtered;
          input_filtered(8) <= in8_filtered;
--          input_filtered(9) <= in9_filtered;
--          input_filtered(10) <= in10_filtered;

		  input_filtered(0) <= input_filtered0_temp;
		  input_filtered(4) <= input_filtered4_temp;
		  
          intr_input_reg(0) <= intr_in0;
          intr_input_reg(1) <= intr_in1;
          intr_input_reg(2) <= intr_in2;
          intr_input_reg(3) <= intr_in3;
          intr_input_reg(4) <= intr_in4;
          intr_input_reg(5) <= intr_in5;
          intr_input_reg(6) <= intr_in6;
          intr_input_reg(7) <= intr_in7;
          intr_input_reg(8) <= intr_in8;
--          intr_input_reg(9) <= intr_in9;
--          intr_input_reg(10) <= intr_in10;

          input_flag_reg(0) <= intr_in0_flag;
          input_flag_reg(1) <= intr_in1_flag;
          input_flag_reg(2) <= intr_in2_flag;
          input_flag_reg(3) <= intr_in3_flag;
          input_flag_reg(4) <= intr_in4_flag;
          input_flag_reg(5) <= intr_in5_flag;
          input_flag_reg(6) <= intr_in6_flag;
          input_flag_reg(7) <= intr_in7_flag;
          input_flag_reg(8) <= intr_in8_flag;
--          input_flag_reg(9) <= intr_in9_flag;
--          input_flag_reg(10) <= intr_in10_flag;

---------------------- Configuration Registers ---------------------

-- Configuration Register 1 
--
-- Controls the input polarity
-- and input debounce filtering for each input signal.

	input_config1_regen <= input_config1_dcd AND not(Nwr);
	
	register1: process (mclk, Nreset)
    BEGIN

	if(Nreset='0') then
        input_config1 <= (others=>'0');
	elsif(rising_edge (mclk)) then
        if (input_config1_regen='1') then
        	input_config1 <= data;
	    end if;
	end if;
    END process register1;

--    in_filter_select10 <= input_config1(31 downto 30);
--    in_filter_select9 <= input_config1(29 downto 28);
    in_filter_select8 <= input_config1(27 downto 26);
    in_filter_select7 <= input_config1(25 downto 24);
    in_filter_select6 <= input_config1(23 downto 22);
    in_filter_select5 <= input_config1(21 downto 20);
    in_filter_select4 <= input_config1(19 downto 18);
    in_filter_select3 <= input_config1(17 downto 16);
    in_filter_select2 <= input_config1(15 downto 14);
    in_filter_select1 <= input_config1(13 downto 12);
    in_filter_select0 <= input_config1(11 downto 10);

    -- The default input polarity is active low.  Entering a "1"
    -- for the invert reg value defines the input as active high.
    -- Inputs will be reported to the software as the filtered
    -- and as active high value at all times, internally.

    in_invreg(8 downto 0) <= input_config1(8 downto 0);
--    in_invreg(10) <= input_config1(9);
	
	-- Need to generate in_invreg(10) from another bit in some reg.
	-- For now, bit 9 controls both 9 & 10 invert sense.
		
---------------------------------------------------------------

-- Configuration Register 2 
--
-- Controls the pulse or level mode of each output and the pulse
-- duration in pulse mode.  This is done by assigning three bits 
-- to each of the six general purpose outputs.  
--
-- For the general purpose outputs the three-bit control definition
-- is:
--
--  OUTPUT TYPE
--    bit(n+2)  bit(n+1)  bit(n)  Pulse Width
--    1=PULSE        1    1       40 msec
--    0=NO PULSE     1    0       10 msec
--                   0    1        5 msec
--                   0    0        5 usec
--

	output_config2_regen <= output_config2_dcd AND not(Nwr);
	
	load_output_config2: process (mclk, Nreset)
    BEGIN

	if(Nreset='0') then
        output_config2 <= (others=>'0');
	elsif(rising_edge (mclk)) then
        if (output_config2_regen='1') then
        	output_config2 <= data;
	    end if;
	end if;
    END process load_output_config2;
	
	output_active <= output_config2(31);
	
    gatemode_a <= output_config2(30 downto 28);
    gatemode_b <= output_config2(27 downto 25);

--    pulse_mode_8  <= output_config2(23);			-- output 8 controlled same as output 7;
--    pulse_width_8 <= output_config2(22 downto 21); -- not enough bits for independent control.

    pulse_mode_7  <= output_config2(23);
    pulse_width_7 <= output_config2(22 downto 21);

    pulse_mode_6  <= output_config2(20);
    pulse_width_6 <= output_config2(19 downto 18);

    pulse_mode_5  <= output_config2(17);
    pulse_width_5 <= output_config2(16 downto 15);

    pulse_mode_4  <= output_config2(14);
    pulse_width_4 <= output_config2(13 downto 12);

    pulse_mode_3  <= output_config2(11);
    pulse_width_3 <= output_config2(10 downto 9);

    pulse_mode_2  <= output_config2(8);
    pulse_width_2 <= output_config2(7 downto 6);

    pulse_mode_1  <= output_config2(5);
    pulse_width_1 <= output_config2(4 downto 3);

    pulse_mode_0  <= output_config2(2);
    pulse_width_0 <= output_config2(1 downto 0);

---------------------------------------------------------------

-- Configuration Register 3 
--
-- Controls the source of each output
-- signal.  The sources include a software controlled bit, which
-- may be written by software due one of several conditions occurring.
-- Also, other hardware sources can be selected, such as print image
-- completion.
--
-- In addition, this register controls the enable for each of the
-- input interrupts.  
--
-- The configuration bits are defined here.
--
-- Each interrupt enable bit is set to a '1' to enable and '0' to disable
-- that interrupt.
--
-- intr_enable(9 downto 0) <= config3(27 downto 18)
--
-- SOURCE          bit(n+2)  bit(n+1)  bit(n)
-- 
-- Software-controlled   1      0       0
-- Image Complete, hd.1  0      0       0
-- Print Ready, hd. 1    0      0       1
-- Image Complete, hd.2  0      1       0
-- Print Ready, hd. 2    0      1       1

-- Now that we only control a single head, we can eliminate the middle
-- column in the above table.  Two bits per output control the 
-- source select (column 1 & 3 above).

	outsrc_config3_regen <= outsrc_config3_dcd AND not(Nwr);
	
	register3: process (mclk, Nreset)
    BEGIN

	if(Nreset='0') then
        outsrc_config3 <= (others=>'0');
	elsif(rising_edge (mclk)) then
        if (outsrc_config3_regen='1') then
        	outsrc_config3 <= data;
	    end if;
	end if;
    END process register3;


--    two_edge_enable3 <= outsrc_config3(30);
--    two_edge_enable1 <= outsrc_config3(29);

--    intr_in10_enable <= outsrc_config3(28);
--    intr_in9_enable <= outsrc_config3(27);
    intr_in8_enable <= outsrc_config3(26);
    intr_in7_enable <= outsrc_config3(25);
    intr_in6_enable <= outsrc_config3(24);
    intr_in5_enable <= outsrc_config3(23);
    intr_in4_enable <= outsrc_config3(22);
    intr_in3_enable <= outsrc_config3(21);
    intr_in2_enable <= outsrc_config3(20);
    intr_in1_enable <= outsrc_config3(19);
    intr_in0_enable <= outsrc_config3(18);

 --   src_config8 <= outsrc_config3(17 downto 16);
    src_config7 <= outsrc_config3(15 downto 14);
    src_config6 <= outsrc_config3(13 downto 12);
    src_config5 <= outsrc_config3(11 downto 10);
    src_config4 <= outsrc_config3(9 downto 8);
    src_config3 <= outsrc_config3(7 downto 6);
    src_config2 <= outsrc_config3(5 downto 4);
    src_config1 <= outsrc_config3(3 downto 2);
    src_config0 <= outsrc_config3(1 downto 0);

    -- modified source config regs. used for single head version;
    -- no need for extra mux range.  Bit definition satisfied
    -- using only 1st and 3rd bits.  Also, wired 11 choice to
    -- same as 10; i.e. software controlled bit.

--    mod_src_config8 <= outsrc_config3(17) & outsrc_config3(16);
--    same modulation source for inputs 7 and 8 due to limited reg. bits
--    mod_src_config8 <= outsrc_config3(15) & outsrc_config3(14);
    mod_src_config7 <= outsrc_config3(15) & outsrc_config3(14);
    mod_src_config6 <= outsrc_config3(13) & outsrc_config3(12);
    mod_src_config5 <= outsrc_config3(11) & outsrc_config3(10);
    mod_src_config4 <= outsrc_config3(9) & outsrc_config3(8);
    mod_src_config3 <= outsrc_config3(7) & outsrc_config3(6);
    mod_src_config2 <= outsrc_config3(5) & outsrc_config3(4);
    mod_src_config1 <= outsrc_config3(3) & outsrc_config3(2);
    mod_src_config0 <= outsrc_config3(1) & outsrc_config3(0);


---------------------------------------------------------------

-- Configuration Register 4 
--
-- Controls the software-controlled output bits.  Currently, this
-- register only latches the eight least significant bits.  A 
-- separate address was defined for this so as to avoid the need
-- for software to mix configuration data with output data.
--
-- For the tri-color alert light, the two-bit control definition is:
--
-- OUTPUT STATE     bit(n+1)  bit(n)
--
-- Flashing, 2 per sec.  1    1
-- Flashing, 1 per sec.  1    0
-- Active Low (ON)       0    1
-- Active Low (OFF)      0    0
	
	
	outctrl_config4_regen <= outctrl_config4_dcd AND not(Nwr);
	
	register4: process (mclk, Nreset)
    BEGIN

	if(Nreset='0') then
       	output_data <= (others=>'0');
	    alert_data_siren <= (others=>'0');
	    alert_data_red <= (others=>'0');
	    alert_data_yel <= (others=>'0');
	    alert_data_grn <= (others=>'0');
	elsif(rising_edge (mclk)) then
        if (outctrl_config4_regen='1') then
		    alert_data_siren <= data(27 downto 26);
		    alert_data_red <= data(25 downto 24);
		    alert_data_yel <= data(21 downto 20);
		    alert_data_grn <= data(17 downto 16);
	    end if;
        if (outctrl_config4_regen='1') then
        	output_data <= data(7 downto 0); -- output_data bits written here
        else -- if the output_data was set to a '1' and this is pulse mode,
			 -- then reset output_data to a '0' on the next clock. This permits 
			 -- software to treat the outputs as rising edge sensitive controlled 
			 -- outputs.
            if(output_data(0)='1' AND pulse_mode_0 ='1') then 
                    output_data(0)<='0';
            end if;
            if(output_data(1)='1' AND pulse_mode_1 ='1') then 
                    output_data(1)<='0';
            end if;
            if(output_data(2)='1' AND pulse_mode_2 ='1') then 
                    output_data(2)<='0';
            end if;
            if(output_data(3)='1' AND pulse_mode_3 ='1') then 
                    output_data(3)<='0';
            end if;
            if(output_data(4)='1' AND pulse_mode_4 ='1') then 
                    output_data(4)<='0';
            end if;
            if(output_data(5)='1' AND pulse_mode_5 ='1') then 
                    output_data(5)<='0';
            end if;
            if(output_data(6)='1' AND pulse_mode_6 ='1') then 
                    output_data(6)<='0';
            end if;
            if(output_data(7)='1' AND pulse_mode_7 ='1') then 
                    output_data(7)<='0';
            end if;
--            if(output_data(8)='1' AND pulse_mode_8 ='1') then 
--                    output_data(8)<='0';
--            end if;
	  end if;
      end if;
    END process register4;

	
---------------- Select Output Pulse Timer Clock ---------------

    pulse_tick0: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
        pulse_width_0, pulse_choice0);

    pulse_tick1: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
        pulse_width_1, pulse_choice1);

    pulse_tick2: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
        pulse_width_2, pulse_choice2);

    pulse_tick3: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
        pulse_width_3, pulse_choice3);

    pulse_tick4: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
        pulse_width_4, pulse_choice4);

    pulse_tick5: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
        pulse_width_5, pulse_choice5);

    pulse_tick6: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
        pulse_width_6, pulse_choice6);

    pulse_tick7: selector_4 port map(mclk, Nreset, high, 
        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
        pulse_width_7, pulse_choice7);

--    pulse_tick8: selector_4 port map(mclk, Nreset, high, 
--        clk1mh_tick, clk2_9kh_tick, clk1_45kh_tick, clk362hz_tick,
--        pulse_width_8, pulse_choice8);


---------------- Select Output Source --------------------

-- Modified least significant select bit so that software controlled
-- pulse output doesn't need to be set back to zero for each pulse.
-- The write of a one to the appropriate bit always commands the pulse.

    out_select0: selector_4 port map(mclk, Nreset, high,
        image_done1, print_enable1, output_data(0), output_data(0),
        mod_src_config0, out_choice0);

    out_select1: selector_4 port map(mclk, Nreset, high, 
        image_done1, print_enable1, output_data(1), output_data(1),
        mod_src_config1, out_choice1);

    out_select2: selector_4 port map(mclk, Nreset, high, 
        image_done1, print_enable1, output_data(2), output_data(2),
        mod_src_config2, out_choice2);

    out_select3: selector_4 port map(mclk, Nreset, high, 
        image_done1, print_enable1, output_data(3), output_data(3),
        mod_src_config3, out_choice3);

    out_select4: selector_4 port map(mclk, Nreset, high, 
        image_done1, print_enable1, output_data(4), output_data(4),
        mod_src_config4, out_choice4);

    out_select5: selector_4 port map(mclk, Nreset, high, 
        image_done1, print_enable1, output_data(5), output_data(5),
        mod_src_config5, out_choice5);

    out_select6: selector_4 port map(mclk, Nreset, high, 
        image_done1, print_enable1, output_data(6), output_data(6),
        mod_src_config6, out_choice6);

    out_select7: selector_4 port map(mclk, Nreset, high, 
        image_done1, print_enable1, output_data(7), output_data(7),
        mod_src_config7, out_choice7);

--    out_select8: selector_4 port map(mclk, Nreset, high, 
--        image_done1, print_enable1, output_data(8), output_data(8),
--        mod_src_config8, out_choice8);



---------------- Generate Output Edge Tick --------------------

    -- Allow pulse out unless image done selected; then only if
    -- print is enabled.  This prevents glitches during software
    -- selection, unless print is enabled when changed.

    enabletick0 <= '1' when(output_active='1' AND (print_enable1='1' 
				OR mod_src_config0(1)='1' OR mod_src_config0(0)='1')) else '0';
    enabletick1 <= '1' when(output_active='1' AND (print_enable1='1' 
				OR mod_src_config1(1)='1' OR mod_src_config1(0)='1')) else '0';
    enabletick2 <= '1' when(output_active='1' AND (print_enable1='1' 
				OR mod_src_config2(1)='1' OR mod_src_config2(0)='1')) else '0';
    enabletick3 <= '1' when(output_active='1' AND (print_enable1='1' 
				OR mod_src_config3(1)='1' OR mod_src_config3(0)='1')) else '0';
    enabletick4 <= '1' when(output_active='1' AND (print_enable1='1' 
				OR mod_src_config4(1)='1' OR mod_src_config4(0)='1')) else '0';
    enabletick5 <= '1' when(output_active='1' AND (print_enable1='1' 
				OR mod_src_config5(1)='1' OR mod_src_config5(0)='1')) else '0';
    enabletick6 <= '1' when(output_active='1' AND (print_enable1='1' 
				OR mod_src_config6(1)='1' OR mod_src_config6(0)='1')) else '0';
    enabletick7 <= '1' when(output_active='1' AND (print_enable1='1' 
				OR mod_src_config7(1)='1' OR mod_src_config7(0)='1')) else '0';
--    enabletick8 <= '1' when(output_active='1' AND (print_enable1='1' 
--				OR mod_src_config8(1)='1' OR mod_src_config8(0)='1')) else '0';

	edgeout0: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        out_choice_tick0  <= '0';
        out_choice_del0 <= '0';
	elsif(rising_edge (mclk)) then
        out_choice_del0  <= out_choice0;

		-- mux control may be setting a new source 
		-- when outsrc_config3_regen='1'; this would otherwise 
		--cause a "glitch" if the new source were active. 
		-- Therefore, inhibit tick during mux selection.

        if(out_choice0='1' AND out_choice_del0='0' 
            AND outsrc_config3_regen='0' AND enabletick0='1') then
            out_choice_tick0 <= '1';
        else
            out_choice_tick0 <= '0';
	    end if;
	end if;
    END process edgeout0;

	edgeout1: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        out_choice_tick1  <= '0';
        out_choice_del1 <= '0';
	elsif(rising_edge (mclk)) then
        out_choice_del1  <= out_choice1;

		-- mux control may be selecting a new source 
		-- when outsrc_config3_regen='1'; this would otherwise 
		--cause a "glitch" if the new source were active. 
		-- Therefore, inhibit tick during mux selection.

        if(out_choice1='1' AND out_choice_del1='0'
            AND outsrc_config3_regen='0' AND enabletick1='1') then
            out_choice_tick1 <= '1';
        else
            out_choice_tick1 <= '0';
	    end if;
	end if;
    END process edgeout1;

	edgeout2: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        out_choice_tick2  <= '0';
        out_choice_del2 <= '0';
	elsif(rising_edge (mclk)) then
        out_choice_del2  <= out_choice2;

		-- mux control may be selecting a new source 
		-- when outsrc_config3_regen='1'; this would otherwise 
		--cause a "glitch" if the new source were active. 
		-- Therefore, inhibit tick during mux selection.

        if(out_choice2='1' AND out_choice_del2='0' 
            AND outsrc_config3_regen='0' AND enabletick2='1') then
            out_choice_tick2 <= '1';
        else
            out_choice_tick2 <= '0';
	    end if;
	end if;
    END process edgeout2;

	edgeout3: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        out_choice_tick3  <= '0';
        out_choice_del3 <= '0';
	elsif(rising_edge (mclk)) then
        out_choice_del3  <= out_choice3;

		-- mux control may be selecting a new source 
		-- when outsrc_config3_regen='1'; this would otherwise 
		--cause a "glitch" if the new source were active. 
		-- Therefore, inhibit tick during mux selection.

        if(out_choice3='1' AND out_choice_del3='0' 
            AND outsrc_config3_regen='0' AND enabletick3='1') then
            out_choice_tick3 <= '1';
        else
            out_choice_tick3 <= '0';
	    end if;
	end if;
    END process edgeout3;

	edgeout4: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        out_choice_tick4  <= '0';
        out_choice_del4 <= '0';
	elsif(rising_edge (mclk)) then
        out_choice_del4  <= out_choice4;

		-- mux control may be selecting a new source 
		-- when outsrc_config3_regen='1'; this would otherwise 
		--cause a "glitch" if the new source were active. 
		-- Therefore, inhibit tick during mux selection.

        if(out_choice4='1' AND out_choice_del4='0' 
            AND outsrc_config3_regen='0' AND enabletick4='1') then
            out_choice_tick4 <= '1';
        else
            out_choice_tick4 <= '0';
	    end if;
	end if;
    END process edgeout4;

	edgeout5: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        out_choice_tick5  <= '0';
        out_choice_del5 <= '0';
	elsif(rising_edge (mclk)) then
        out_choice_del5  <= out_choice5;

		-- mux control may be selecting a new source 
		-- when outsrc_config3_regen='1'; this would otherwise 
		--cause a "glitch" if the new source were active. 
		-- Therefore, inhibit tick during mux selection.

        if(out_choice5='1' AND out_choice_del5='0' 
            AND outsrc_config3_regen='0' AND enabletick5='1') then
            out_choice_tick5 <= '1';
        else
            out_choice_tick5 <= '0';
	    end if;
	end if;
    END process edgeout5;

	edgeout6: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        out_choice_tick6  <= '0';
        out_choice_del6 <= '0';
	elsif(rising_edge (mclk)) then
        out_choice_del6  <= out_choice6;

		-- mux control may be selecting a new source 
		-- when outsrc_config3_regen='1'; this would otherwise 
		--cause a "glitch" if the new source were active. 
		-- Therefore, inhibit tick during mux selection.

        if(out_choice6='1' AND out_choice_del6='0' 
            AND outsrc_config3_regen='0' AND enabletick6='1') then
            out_choice_tick6 <= '1';
        else
            out_choice_tick6 <= '0';
	    end if;
	end if;
    END process edgeout6;

	edgeout7: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        out_choice_tick7  <= '0';
        out_choice_del7 <= '0';
	elsif(rising_edge (mclk)) then
        out_choice_del7  <= out_choice7;

		-- mux control may be selecting a new source 
		-- when outsrc_config3_regen='1'; this would otherwise 
		--cause a "glitch" if the new source were active. 
		-- Therefore, inhibit tick during mux selection.

        if(out_choice7='1' AND out_choice_del7='0' 
            AND outsrc_config3_regen='0' AND enabletick7='1') then
            out_choice_tick7 <= '1';
        else
            out_choice_tick7 <= '0';
	    end if;
	end if;
    END process edgeout7;

--	edgeout8: process (mclk, Nreset)
--    BEGIN
--    if (Nreset='0') then
--        out_choice_tick8  <= '0';
--        out_choice_del8 <= '0';
--	elsif(rising_edge (mclk)) then
--        out_choice_del8  <= out_choice8;
--
--		-- mux control may be selecting a new source 
--		-- when outsrc_config3_regen='1'; this would otherwise 
--		--cause a "glitch" if the new source were active. 
--		-- Therefore, inhibit tick during mux selection.
--
--        if(out_choice8='1' AND out_choice_del8='0' 
--            AND outsrc_config3_regen='0' AND enabletick8='1') then
--            out_choice_tick8 <= '1';
--        else
--            out_choice_tick8 <= '0';
--	    end if;
--	end if;
--    END process edgeout8;


------------------ Generate Output Pulse ----------------------
-- pulse_rt_1ms is a 4 bit counter-based retriggerable one-shot

    pulseout0: pulse_rt_1ms port map (
        mclk, Nreset, pulse_choice0, out_choice_tick0, pulse_out0);

    pulseout1: pulse_rt_1ms port map (
        mclk, Nreset, pulse_choice1, out_choice_tick1, pulse_out1);

    pulseout2: pulse_rt_1ms port map (
        mclk, Nreset, pulse_choice2, out_choice_tick2, pulse_out2);

    pulseout3: pulse_rt_1ms port map (
        mclk, Nreset, pulse_choice3, out_choice_tick3, pulse_out3);

    pulseout4: pulse_rt_1ms port map (
        mclk, Nreset, pulse_choice4, out_choice_tick4, pulse_out4);

    pulseout5: pulse_rt_1ms port map (
        mclk, Nreset, pulse_choice5, out_choice_tick5, pulse_out5);
		
    pulseout6: pulse_rt_1ms port map (
        mclk, Nreset, pulse_choice6, out_choice_tick6, pulse_out6);

    pulseout7: pulse_rt_1ms port map (
        mclk, Nreset, pulse_choice7, out_choice_tick7, pulse_out7);

--    pulseout8: pulse_rt_1ms port map (
--        mclk, Nreset, pulse_choice8, out_choice_tick8, pulse_out8);
		
	level_out0 <= out_choice0;
	level_out1 <= out_choice1;
	level_out2 <= out_choice2;
	level_out3 <= out_choice3;
	level_out4 <= out_choice4;
	level_out5 <= out_choice5;
	level_out6 <= out_choice6;
	level_out7 <= out_choice7;
--	level_out8 <= out_choice8;


------------------- OUTPUT GATING LOGIC ---------------------

-- General inputs 0 and 1 are opto-isolated; 
-- inputs 2 through 9 are logic referenced.
-- Outputs 0 and 1 are opto-isolated, outputs 2 thru 5 are logic referenced.

--   gatemode_a(1)   gatemode_a(0)

--      0               0           Gate_A disabled, output active
--      0               1           Gate_A disabled, output active
--      1               0           Gate_A enabled, using logic input 4
--      1               1           Gate_A enabled, using isolated input 0

--   gatemode_a(2) -- UNUSED - GATE A ALWAYS APPLIED TO OUTPUT 0
--      0           Apply gate A to output 2
--      1           Apply gate A to output 0

-- Let the external gate be defined as active to inhibit;
-- inactive to allow normal signal output to pass.

--   gatemode_b(1)   gatemode_b(0)

--      0               0           Gate_B disabled, output active
--      0               1           Gate_B disabled, output active
--      1               0           Gate_B enabled, using logic input 4
--      1               1           Gate_B enabled, using isolated input 0

--   gatemode_b(2) -- UNUSED - GATE B ALWAYS APPLIED TO OUTPUT 2
--      0           Apply gate B to output 2
--      1           Apply gate B to output 0

-- Let the external gate be defined as active to inhibit;
-- inactive to allow normal signal output to pass.

--	input_filtered0_temp
--	input_filtered4_temp


    gate_mux_a : selector_4 
    PORT MAP(mclk, Nreset, high, 
        high, high, input_filtered4_temp, input_filtered0_temp,
        gatemode_a(1 downto 0), gate_enable_A);

    gate_mux_b : selector_4 
    PORT MAP(mclk, Nreset, high, 
        high, high, input_filtered4_temp, input_filtered0_temp,
        gatemode_b(1 downto 0), gate_enable_B);


------------------ Select Output Pulse Type --------------------

    out_enable0 <= output_active AND gate_enable_A;
    out_enable1 <= output_active;
    out_enable2 <= output_active AND gate_enable_B;
    out_enable3 <= output_active;
    out_enable4 <= output_active;
    out_enable5 <= output_active;
    out_enable6 <= output_active;
    out_enable7 <= output_active;
--    out_enable8 <= output_active;


    type_select0 : selector_2 port map(mclk, Nreset, out_enable0, 
        level_out0, pulse_out0, pulse_mode_0,
		gen_out0);

        Ngen_out(0) <= not(gen_out0);

    type_select1 : selector_2 port map(mclk, Nreset, out_enable1, 
        level_out1, pulse_out1, pulse_mode_1,
		gen_out1);

        Ngen_out(1) <= not(gen_out1);

    type_select2 : selector_2 port map(mclk, Nreset, out_enable2, 
        level_out2, pulse_out2, pulse_mode_2,
		gen_out2);

        Ngen_out(2) <= not(gen_out2);

    type_select3 : selector_2 port map(mclk, Nreset, out_enable3, 
        level_out3, pulse_out3, pulse_mode_3,
		gen_out3);

        Ngen_out(3) <= not(gen_out3);

    type_select4 : selector_2 port map(mclk, Nreset, out_enable4, 
        level_out4, pulse_out4, pulse_mode_4,
		gen_out4);

        Ngen_out(4) <= not(gen_out4);

    type_select5 : selector_2 port map(mclk, Nreset, out_enable5, 
        level_out5, pulse_out5, pulse_mode_5,
		gen_out5);

        Ngen_out(5) <= not(gen_out5);

    type_select6 : selector_2 port map(mclk, Nreset, out_enable6, 
        level_out6, pulse_out6, pulse_mode_6,
		gen_out6);

        Ngen_out(6) <= not(gen_out6);

    type_select7 : selector_2 port map(mclk, Nreset, out_enable7, 
        level_out7, pulse_out7, pulse_mode_7,
		gen_out7);

        Ngen_out(7) <= not(gen_out7);

--    type_select8 : selector_2 port map(mclk, Nreset, out_enable8, 
--        level_out8, pulse_out8, pulse_mode_8,
--		gen_out8);
--
--        Ngen_out(8) <= not(gen_out8);


-- OUTPUT STATE     bit(n+1)  bit(n)
--
-- Flashing, 2 per sec.  1    1
-- Flashing, 1 per sec.  1    0
-- Active Low (ON)       0    1
-- Active Low (OFF)      0    0

	flash_timing: process (mclk, Nreset)
    BEGIN
    if (Nreset='0') then
        flash_count <= (others=>'0');
		half_sec_toggle <= '0';
		qtr_sec_toggle <= '0';
	elsif(rising_edge (mclk)) then
        if(clk181hz_tick='1') then
			if(flash_count="101101") then -- count of 45
				flash_count <= (others =>'0');
				qtr_sec_toggle <= not(qtr_sec_toggle);
				if(qtr_sec_toggle='1') then
					half_sec_toggle <= not(half_sec_toggle);
				end if;
			else
            	flash_count <= flash_count + 1;
			end if;
	    end if;
	end if;
    END process flash_timing;

	flash_1sec <= half_sec_toggle;
	flash_half_sec <= qtr_sec_toggle;

    flashmuxsiren: selector_4 port map(mclk, Nreset, output_active, 
        low, high, flash_1sec, flash_half_sec,
        alert_data_siren, siren);

	Nsiren <= not(siren);		

    flashmuxred: selector_4 port map(mclk, Nreset, output_active, 
        low, high, flash_1sec, flash_half_sec,
        alert_data_red, tri_red);

	Ntri_red <= not(tri_red);		

    flashmuxyel: selector_4 port map(mclk, Nreset, output_active, 
        low, high, flash_1sec, flash_half_sec,
        alert_data_yel, tri_yel);
		
	Ntri_yel <= not(tri_yel);		

    flashmuxgrn: selector_4 port map(mclk, Nreset, output_active, 
        low, high, flash_1sec, flash_half_sec,
        alert_data_grn, tri_grn);
		
	Ntri_grn <= not(tri_grn);		

END archiologic10;

